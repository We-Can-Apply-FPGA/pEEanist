��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��`Ղ���0<a6B��(I�izr��6����,��_��M�:��&�PH���da[��a���V��z��#��bV�#~Z�T�����K���]��v�Ÿ����e�Ǐ�U�F����XPd�}�4T���|�������~"�l�A�]^^R�2.���1ח��:bZ����Q�E/4:�He��"`�XM���xǑ�/��(^H��v6�j��2��F�爴���9�2��y��\�Ob�w��Ne`ӷSK�z�41B���٩d#�*����]�o�܇u1@bMJ�L��2��]u�:#�!̘��*|Q���24����k�)a+��upg�9"�bl@Α�z�y,���q4ꊙ����A;�z�>�X�ruI�7���<�A���s�A{�I�6�6�iV\F�E��o�E3Ef6g��1[x\��[I��Ai��&hSڡ�"fIw>v6HXVp�c�_PD�^�oD����H���].���uH�]�.�
���t��zP\��@�C&��
	��U�E�jv��j�ɱ�Aoj���#4����fv֜��}wVmV�|u��9�.�O����`r�h�D
�k��r���H����?h�H�*)�VyA���\���=4dK��y�����B4��2�mm#��G��:j������T�0N���yt&1�yk���� ���L�mP�A��ޠy`�}�ESz�z|�F�m�u��*Ǫ@@�w �zp�	�E�]�R��{�=y�eM0���3۩�s�L,�C+k_��N�����.�	�+�v�������G/"<��$N���=0�J����XmXV�=��֬U��)}ꁜ�oL����f׌�'r�e΢���W��ߞ�797I�+�Fl�ԓ*��@�M
]�h�,���r8^P�E	��"'�L
ӏ�}�DYKuB�׸'�dٜ�������5 ���g��[Ԫ'?��� ��P6�W�����.����
�vNaH�g%�o,�k׉�j�vMw��T;�@��h�b��R�ՊBA���&U:����eu�t-b{�m~;$��A%^�����m�E�(�w>]�W�����͛Y�=�~��>�予b
�� fe.dfi�3�֮K~I�r�U�(��g�p��;dk�v�³��X%fP�ڠ�>�.)��\�zf��E���lQ�l��s����9G�x�_�_��~����1A_q�d�!�sV#`Nr�Y-�I�M.={�����[]�`Z͖ߌe0*pK�1,�NK�ϱ�h��t�tL�WV���4(7�1vx5t�Ez2A��fC�&:��m�.��}���+��Tdm�cg�Dƺ�S�._9���3�w�g[_�>w ��g�wY�Z۞Կ�Q]1P�,�g���Fѡ��Ħ���UH�x���A�霟<öo�2���Ldl��M6��FְC;Vd0g��"ɡ�oY��%v�	�ĸo�*������?FH_�S���f�q���g?�a�͚G�A�Q�>C	]���=���F����G��"�aИ<'��76i�4L[A�3u��]����G/�ň��Ue�w_�?"$ú�s�i?G¨�]'��e�67��x�����(�32ж��vr?#}J������]�o�}޶��K`����B��g�/�ݒ|V�m�nm�g���懁{&���[|�EY����V��3��U��/�"�0��������"{;��h:f���ij������txB��o��=��|�F�����a�h�w06Ad����S`�p ����N0��:�u��f���le���bu��7XÁ���	��A�C�����%�?�坈�W8��=z�]���3���$-{}�jE�	�Wn�ыɔ|��I	��!M��9g������ɠ�Quz�:kk����G^�4EV�s.��"�m[�Y���b��WWc�d�θ��I����m��bC7�X^�|k"��'?|,Kh��a?=����=㬬k��{J���b��_J�S� �%�mMU�+6m��B�"��kᖁ�S,+�W�D�Er]&+K]�x-�At����^&��U���d閖��g//��d����h�u���Ý�����i��Б"*��(^=(��V�!%6������HXs�*�_��S�����$���{x�ˤ���;�L"Bo���Շ�g��D����ڊ��ix��a�*0C��	AnR2�M�0v<zX5f��8��s1{U����m��p7)<���x��<���;��P�/$�n����oH�#�VD�V��hÃ�cY�����f���y��[��؃8�F:�4��TC��C �VN4��.%�����? ����f�ŵ�΂L[/)�7R}T��豕鸝U��n0[�,'$�����U֥�1J���t]K�ʷ�t�pvР��?.�'�Dgm�����_������8�]x�!Ņm�0K�/TDS?ڦR�ʀL_�%J�~SV��q�7��{���џ���AO��pBc���C�"�K�����G��d��K��/��n��X˹�$�E���0 N�8Ԭ[�c�*� :a�c�|����q��<���PmW��`y���z��y���Q�u
�sq�0'�!��녳�L��`�fMj��ʰC|V�4S{#�eH�(�QJM5C�;��4:�e��i|y��A����62��F\��%⛡w�WG3|w�p��S�Ґ�X�j2q�5�"�wҺ���4`���־����Q��̪ܺZ�XO����Y*Z��E!�������̚M��N�S��k;l1�tO�V�������P������m=���Y�� *C�Ƙ�����m-�W�  r�{7���<B~��)���k�Jq�aK��"~2`H���������a@�,a�XK�I�
�~E�,P1^���Z.�Ga�Q��䋝�B�w�w`Y>X?��Y����s9�T����C.e�#����.���&@7���O�U�Y����7�0`>�<��<!��y�Y����E3��E��r��<x���Aۈ��,Q��GpB{"�u�&��S�R�o򧼾X�3��R�\*��S�~���V�ls���U��=��P�`�=~��eK(�g�݃�Q�=ZLPY�\�W])�*���:T�;��s	��t`�ϮA�0��k���2�i)ft=Q�#�����z�'ԍ�*��NO��6m�m(���f��]B�Ɉy=!���||
��U��͸�M�H��+�9�]�𛼁�UU/�5@�$�ʣ���pF;�u�͝~��
16�Z�>��#��@���^5!�q�K��k~Y�9P[Ł�A�ԨŦK{�܃���X���3o2��֎���TT69ݒIJۦ�)2�V��b]����-�����}6�f�3�i�����Xf����m�?���Q��F[Re�T����.~�vE�,�<*aK��������Rt#��N����V�y?����x�À��-��O��fRU�N�%8�����e������B��q*��_��8�-�.nR�v��B�B��}����	S�z�c�)">cG7��b)!���Q��,r^/ʢ�^��gV������/�����
���7��������)�R�BDA�+}�V`N<9�@���B;����a����Ta��\����w�S0 3�4�V?��ߖ1�V�Z��U�:���Y)!@=xظ0I�E]���u�Bd��E�3���o��XH��`鋶��}�yga���c\����g.�T5�8Q9��%	�*��}�S�� �`�Y�p(�d�M�����qM:|
�/n��!�������5�u�5,p t��7������(ܟ�?���?zeH���"������pm�bׄ��Rx�R�� M�*�O�Umwa�J�|�9Ɇ?QC�ء޿
'M�� 62C�Q^��ɤ5�����bM� Z^��D�AJ�0���_��������=4��s��M�a���R��lX4��ށn��	�q��m�����@�x�h��Q���\?޴�yn�ec0��.�[7܆������� Ηun��G4޻YQ�i�yo�R%����
R_�|� �U ��DXT�Ħ��_p�U4�9��e���2��q&�.qx���yGat�z��r7��k����AO<��օ�OY�
0�#!p�^@d�Q5�ףq*�J(r��ю}�(u���H\Z�=��A�O�T� ;�ps�b#MXra��o��s8�e��Wp�G)�ރ�i�{`�r���,���%W�ɶ)���Lv|�脲�JUҹ׆��?-\T���ǆ
�"E<��Q'�+;O�%�k2��i4)��6�Ҷ+�,�)�x�5���	B�^}����&�&���Z3�L�,��.�DQjӒc-�^��%�i2��� Ue~�$�/���0����i;T��P����%��ɠ͏��%��{�^ �U���6Q���;���T�7��n�����w�G��D���L���Z�n�>KA(4��aral	�����`\c�}�?�"�LaL�VQg(��SnW�!S�s�ba;�,?<���g$�hD�B��	�'Rg����ɶ�J��a����Q:\'�.>�n柝L��k���,Z�<�rZ��k�X��T�m��=���yj9G�
{�<Ө�
���V�ƍ���ہ,�	2��7����k9?J)��r7SY#�Ս2M�N�c��/�2ON��9klЏ�
2�٧��c����h�)YQ�]�RlO�r�1g��,�S���h�.�=���E�{�Y��Yci�n��I,gj½�p�� ��譝<�J�X��}�Y�6<�����ݥA�:�D���@�z��?۱0}Awq�G��E"��}L���H�PVE�^�f���Ͱ?��<���h���>��W�������Y��ď�MA�&��M.�b�)����oXO�X���pbk�o-�l�0��=���D���>}n�l�M�~�
"}H�w&󅢆w/��~#� ���/_Q<���ԛ�f�^���(>�	p���-��.�Q��f��~�\+0p��eW�Ț��un'd���.�+�@�0�g����<� �����h)���Bo��VIې�E Y��Amh.k���!��ƿ"�R�$3���I�#S+��f���e(��U�����������GJbS�I�2j.(޾��8�9�w�Rv���"P���a��&��k�����2j7�S�^IB��HV|�b�����eϒ�8a ��2犆����M܇C�V'�#�br������@�%1�=����H�D���@�+�$^l��x!���/��		�����d ��Pa���s�o�[98q�"i���8���Ⱥ\~�Xr
��/�Д�=�Z)OtNI#�J=n���C���v�/(��H�����۽-J-�([0q	1@l���ҿ*[|&(�{����Ã��*�?B1�Կ�d��P�m1��h��PM�dQv��m	X��V�=�p��,�Þ�����f%���N谝[U� �igvN�����[i�M��'3���i�,D4
�Y5��Ҵ��P��A�-��6�e�Ǳ>�|@�6j�K=�$p���V! �D���d^̱��[�]�&+A,!�t~$�m݉n��cM�g.�nt�z��_y��U�*�_[�:QV�<���_��`���Wu�M���x���	Z��  �ӭ��ߨ�	|s%���`ؤZ����9u�NF0ws��*\%��Ý1sp\O��6n��h�M�=�By�Z��z�s'����F9�H�db2�ĸBv�Mړͻ����}P2�.^���������A7��ϣ��Ȃ:8�ßZ3YW!��¤?���4#�+�L���>y_��%���]�`�m^�Y2��k�;��"�v6��!m��wY��vZ���y�\�Px�g#KQ���׉�ğ�eg���R�,ҡ�t8�j�]Q��wN�e��*]3�l$�ˬ�qC����:��7�g7��ؖ2��H�W���=&d5����O^����~A	/=�9r�ws6�dk��`�S�Ά?cZ�w�������3�����a�y|}h�v�4�;�:�6胑tZ��t�N���_k���ڿ8�S��b����Έ��|e(R�+N�~9�DC��X�a�ݕ!Z��|���q�
Ē�g#�ߐ��YD~o��v���}��	�AB��D`��{�H�u��;��k�]���(��c�x,�)�#��Ո��o�>�'��/F�ޙ��m7j_#�=�opW�1���:6!HM�Ӆ�Q��"$6�n�f��ej��a��q{��Y}�*.���5�Z�ȼ��E���� �z�(���~z��#* �M�:��]�������"�;��V�l�����7��[7�R���"�rZ�)4,���̳��t0���
xle/Z��7iu�$t�p�%���m}+�U��Z�H��܁�4S�=�6$b�1���9�o�L��1�i�{i,� �\��F#�Ɋ��:߂�E��= �)��S0��_cx$:a�&FN+�	_�k�E�wR���)��]b�+��r`��V�.4x
H��$uS���ڨ�k���w�TF���-
q�W��k��6#OL訫�Gt���T!��xnL�IkƗ��qQ\��T�k��E�eٱ}��q޽��D��.��Dy��<j���8+3�Mb�-W��u�!{Js���t��US:����7�u&%�V�/�w����N|�m�����Pt�,��;�6�)>)K������9��ύ��{'����QY�����{�Q뽇jڼ��e(�S�1�bi�ŦE��u������s���\=�8c�r�����ia �#��1m�p?����"������Ǳ�
���("\�eH��J�L��
�����#�݃�b!�NC�<6�D\����)�Y�X&[d�r�`9|H��-C���D�;ڣu1��RA�N�o=�lBX����;�v͠��Dd�		���pDXt����X
�IK�Q��n�2�	Of��<{Lӥ�{����c7���& �-k�Bᛵ/�F���F+�F
�M?��W t�;bD|�A	�A:��@ͯ�f�����l�)YCR��}U�`)W%����r���o�V�s�K�s@*��>����Y�,X�K�9.�4���+��OY���6)���C��ǷBea�<u�Ԛ��u���;����5�x�'������QC�{_Mr4���vJ{��X����B��ifqeD	��=�˙�.��&���-n�'{*?rz�@9�UnI1|�W$sv4#�)�ƪ)[�{֙|�Ox���T�A�s���"-j��u�N���1?�n��s W�L���W4��{%.��kp=�J	���Вd��N/l�'J9��-R����1frT�Q��{�Q Ssvh�/8֨aج=�����_^<����VX}��k�(�֌�C�}7;�,�;��\��CR����)�֒ṃ�	�t�4��gp�*{SJ��}"3�؄t�F*p�N�XN����<Mq�����H���7	Ꝯ&n{���83���"K����6-������m1|� L�6��.[]�+֑r�OTu�h[ʕ�=�3cl<!�V<.�A�.@��ہ�O��5Ns�%�Ȥ?սq�U�� ��oP�|�V�z-���O��a�(�l]���9'�9zC��E�v�����Y��iKo�k�T��-tbu5{�:}\��ݝ�j�P�e ��˕ȱ��]e�ߴ�P��*��w`cQ��|XPFd�ĭ�a�
���L��Ƅb���,z�F@�q�ʡ�f�:$`į�K�l�eJo%��#���':𳔹�mY�	b�K���D�X�R�&�|��X��`�݉UT��D�SC3���J��Ѡ'�o��G��}��Y����$^�J��%Ɔಊ�Da%�d�@��=��BE6�=Y��Po��&,r`��H�P���⟼@��($�d��noՋ�4�G7l���*1��*m��=@�����D;`�l�:0J����eM_.�tՀ�]�Ն����k��<$��9��x!ĝ��tr\���-k�T�q���ī����� ���H����F�6xҝb+ro�eZ#����w�7�&�r�2^/�'���eAl%���n�χ�Z�4�_�!'Z(�Pʈ�o�Ǟg��Z� ���/̳e�'���,��At4sc���j�B"�`��(D�&1�b6�<EAv+5�ڝ�Ŭc���`�mS6Q!��Pq�sa�\c[Ƹ�S��it'�x��z��cO�$_��������Ѭ���ܮ,�4�G
�&C�ȟ�$>��>&�G�gY��r�3��0���tұK���\��!� V=j �W�A�륍��yZ�M�� Q�F�b�z�!�q�xL+k��q�<�������j��>d�:i`�������o� ������FzF�i���C�ҠQ���;�V��
$�Z�e�.p����%4��NP��#�n����/2ë[B�P]Ti���6�l^ӪA�B�G4i������P�,~C�%�fZ�a`�F�0 � V%H��j�xV:MP�ij&Mv�+&�|lk��r����K�>BG*ߑ
�������kX�Y=o ��H�^��
�EBK��%��n�R� �_��H�4���-3V]���N#ܕ�2V�I8�Y��Ctn�)'�KY�|%,	��3�X�8X�a�X=���+c��^s-�>�v���C"��/}T̎D��%F�h��]�e�W��s��@�y��{��I6���,��7S�(�!`(��/���I5��O�	���]�6 @�7�l��Ǳ�$SN4�4x9�|&�2����կQVu���(�H)�:󉟅]�3��4�t�p�]v-��3�0��c�M7Z��p)%�@\�]��F1&��1�����A��|ź���d.����6���B��8M����l'��c�g"�	�Ո��ҿ,D;��fx��kJ� i��	ۥaB�	�N��A��h��k$��&YLv�ۡ�հ��tW�?���r����e�.�Įi�N����rǤ$�f,׮�  iGb1Ι�'Ú������
�	��P��?ʔ����{��-׉�Z�䩌�N�0��x��׏}��H5fTٰ(R. Z�pŒ��˓����H�a�����-zCOk�%�0���G����4U�e�()"�	Y�/8@̦��3d���m�"c&�v!�~ˈX�,��I|)���k���f Z��r�mmox��ީd�`�6{�l��x�g��|i[E'��[��}�Q��FG�>�Y�a}�f��{{!�p�ii���~V'z�]��1����Y�/?M��!t��G�C�n!�v��t�2R|{��K��1��QyU��C���`!�2��q��3gC�� �$������_�Z?��o�*���æ�_q,1�db��4�5&�")~h�ay�����%z2�'c"��H�&$*-A���[��=��4c��̳��	�p��q�8^k�[D�*A�1u^"a;h�y��4��Fs-o���x�B	�|c�SK"��!_v���^�΁�å�����iQ���n��95�m�=�2�Xbh��y?��D�7�|��M���d �3�����LF��D����4:�}�L����:��'��=�I�U���\l�Eb��ew�⿦D�4`Ci͈������;��a�������p�W�ܒ3: �+(<�Y�(�K7F��6;\�w�e�D�dsҊ�Җ#獦�1�UAR<R�*LE����{":��A��>ae"#��GP>z2V��j�%�Dؔ�_߳����&鷜��	q@$c��X*e�ro@������4������������#��RO�|ʣ�HN�a�G���u�$���7��
"[�o^�㍱���I�S�8�S^d�b�,�%�a�6�,�������7F(��6�>�.�o�v/#vZr�;r���c]�=0m� D�����$C㑣������Gtx����h�f	!5�c�]�&U`�j��kTJ�}o��v�_8�e���4W�A�,��:1��? �`��і��ɸ8W�70�wR8�gAW	̯�G�a��g"���U�Pc�������E��#kaЋ��eX��jAY*��@�$t$����t������@#�S��T�z�kQR�D�D�)�
q!�y�@1����s[�Z�W!1f2�
v�+�T�&�y�0��}Q����-����;��~�E��Ѧ��e�b���d81�J�T*[	G��	v��TT��א{u��/��AܘFS��u�7�����rP؏K0�4.�6xQԬ���vuVRG反n#Pυs� �C-����G;ra��a=�4�V�ǎ�N$�����n�a����X)H棧m@��\H�؄`Eh����.,�X�ʆ2c���S�0��"��@�Z۵n
�6n9�A���^�y}l7���'�r�=AK�����D�QH�G�K=d<{��Ug QH0��FPqq}q��>��������G��o_U7
zp:"	:n��>�d;�+��{�c�>�e��Jz��z���d3&�y���H*&�`��;�5g�CHt�<��h"�����й��l�n~QE/j�Qx�s�#︭��9����]���n����\= a������D��H��N���3�Ke�5|ZBnz��:�<����GdS�X�`qWC����w�b�#s�r<�9&FXTs,q�!  x�����-?H��c @��<��KdzB�Gڃ��Y`��3�a���S��+��f�؈�W���6R3�^-H��k+��Y����ċ��)I�L�7-t�>����l�~wʈ�P�hå��d�f�
��tYpj��7G.�>��h�����l�>i��kc�Z1>�*�pZ�"�D�*$�/E�2�`~Yul���!�V�����R�AϫU��]F��Ub�m�ԟ},�Ѿ��o��s][�]ؑ�w5H!�\�P�uhbW���n麅���P���h��C��W��TN$��E�I���?R|,��N
��i����7WF���+�t�p�WL$�%I���;�U�"r\��$�r��>��HL����u]�^r*I'�=s%��
Z�4�]�Zk��aX�#R4�z��g��Q�� R4#Eh��F�m^�+�V�Pt^>Fbfg-��r
�H�d�刢@��B\?� B�j�#���78!P?�n�xr/u�CZX���j�ZZj�	���[��b&�pP��Y�S���l5��o��jm�O:���m)�LKN��2{��y+���Ik)�RlN�������� U�{����^��q��p�3�
5B�ʹ�����C��4��M��+���X<%������|��o"�� ͬa�cx"��a^d ����s�'F�G� �	c��l.���G���M�����&�j3?^��@���w �<�j]/o�Ù�������:�pʭ�#�(��PJe���V88��,�l�k3�\t?��Ԝ83�Ǚ>�-�'���1Rd��-�[��(� ����^���ۂ�7t�f�j�HY�w�(�=�eܟ)�v�y	�^�����a�c��O]r���^!���s�<wF}�~��H��[4�2҄d� ��pͣ8������l.�)+"(:m�
<��tĪвU��n�^·�=��S�׻U��U	w�d����UY�8��l׽�̠�$�+@�p���[�z_o�Y,a�4֦Z>���+���Z�u.�T]?6g T�s���cB�?ԕh�~�̨��)C�zH:Vχ/5Y��4�3��1����T.�T�X�	����g@wZ�J�799��^���N������o�(��ºǯ&��=�P&[5�尲Yhe�Aׂ�������r!��}ri�h	g)4��l�Hd5мBs��P���&K���'��y�8��0Uv��7��n9Ő��/}V^o@��Jbq�P!���N-�l�-L@c@������8Q�X��sC��ύWG؛�G���I��G~և�'hl`�ԳuW��>�=��C�Vrʲ�ֶm���)��򆬆�c�Y��E4�z��EC�(���Dn������C�;��__�b�aK'���Z��J"��QT�7��w��?�� �� N147'9?��] ɥ��V��:�ԉ��1	N%��8`q�A���_!�t��2��c�e��G7P�s���u/oC=>'�b���c��v�!Ys��]�N��[w�(����WԕJ���f9W[��=
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i��������쀞L̓"�oܜf�~�5@�g4�5�	�
����,aeH>)�3+,���KԾ�D�X��x���ark��!��H�ҫC��\���!Q{���,�1�Y{�fd�wGP�n-���"����R�j��{��Ҏ쬟�b�Vji��a�a�n��젭Y�?T�K�1����MY�`�4)���Rg�O�C�p���5��la�Dv��F�EC"���L6�ܟo����{H����u{١l�hLk�輎A��m*����x�SN�8�F�S3�k�Q�͟碬��� �� 4L��
T���#YEQDWP\�9�ڛ��ܚV`]������dj��p�ETZ@บ���9�fފ��[�8�o��esO�/�nIӬ�S��k�m�g�7����	���540�m��p�k(<���{n���o	+.aq<P�Y73G��� ���md3�#���g Q/�JI�S��f2H���	�^n�.>��DL�h\������B��A�63�v� j�c��A ��tZ��<q�M٫�œT*��-8u�6d¥�O3�'�bK����ؿ*u~�:Ā�5�����7�KE�f⳨���Hz��qOBd�u@y#q�Q����3���9:ț�N�����V�6!ו��=��I�@$��Z^��'��E��y�*H���[hc���FG;[˙��wmlf�rd$��%E��ob�����,����$���b~�q�#�P�Iw�и� o|����zI�ʂ�Q	~���N-����D&����o��h� bT��6;T�,���� t-u?�0¤��rY�DXA�}�H���:m}c���Q��@{F��!u������
y���l�7MVZ�ߜ��&9�V^I�5���qm���(MtA��P��d�a�Hh��p6�l
�t�L97{�3�|>�R�r���)0�j������N+�cJ3�X�D"T���6>��.�g��$3���f�����p��(M/�,�E'rН?�݈��`�z���Ț��>j������Ȍ�zZ��ɧ%�9Wߺ�2廙׌]��̄��쯨�<�D�'$�Xk`$4��@�V�.� b!�l'j��b	�c���Ge�ő8߫�a �&�^f�J�]��A���8�zt�?��tWzBQ��,�փ�bԢR�����Mp�k���%��g{<%��	�a�m�y��%�j�b��B��S���X}����D2���y�d���<�7�K����V�VO�	j*W�h��3�L��g=%l�?������k#��@�IqU+5m=Y�`���;-�;wϱ/U+���!��:�g�(���~�յ��T� �|KUu���k�*�>�]Ű�q�<Oh cx+UZ�A�xx�+~lN`9��HBJ�~%�?z��:���Qq��|�����)���R�<�?@����	��eKW�y�2���1����n��%&���D��փ��=�U�Sj8��fu.I�<�r���q�e*d^<�=��!#�Ä��ˊ'R�T�$ ��|#���	�VQ�[̡�j�d��M��^j~�5�Mr2���^lo���x�cr�����͍�R�nɑ��\a4�|0�L�Ѧ�'-�tf�\m<t�u�r�?��Y_y�S���&T�� ��4�ʽ�6E\-�P:/�%(��6J���h[Fg
7�#���5����z�$=#�$5����C{�L�e�O�P��~�eS����'��x�r���ܚ����iʵ��0�
�g`���m��m��J������7!e��t�_��kVC(�X1%y��a]���ob�N��^�ݰ&ku�xOo��O�!���o!����8�M^�>0�r�3(S7ꞝ*�篒Pϯ���[�/�@Á��������T�����7M��g�9������iJ-)ƹ�5@�Z[�-��]�T\�o�d��u:}�� �������P�ĆY}�o�{�ci&���ĽC�1]���w3_�� ���*?�c9F?zDb�v�a_HP-�G��2�g����{�3G����u�#�%%5��s���Q���ݭlg��/�Y��q܍����*�|�y�
е��pk������㙐w�V+�i���S���i�V�y<T�O�h����P�� �V#�K�w����g�Dd����uթ�-N6�&oV�2�jŴ4R'���s��<��Lϐ�Q��N�hey����0�!��o��5>�13jw���~!�e�%����ܽ��#�M)P�X��l"P;(J�q� ��.M�1�U5�1(�XY"��t�0t�K�S���/x�AL�hb7�,��p���G��M�k� �Rg�׫��3��@�)������R�ż`&B`3�~xK�n��k��$* >c����{�ɿH<�z� I�:`�N��XJf^�z�MHɲ�먔)�S��a�"J��m2�M�L�G-��+'&6���(S�j���?Zx��;
�B�KԆ�mO5>�8�w�i�3��a�X���.օ�n���<x-v����$"a�V�k���X�o���%X[�f��ϪT#b.�X�"*�I;��͙5�P!���|��]>�2d,�Ub��E��e��o��V��"�'���dpA��\u<�W��!�=�뷜�L��Ž��:ͤGۦ-ZbS��7����<�O�0j{�'���� \��� zX�Y���_�%�(pe~�b�Jr��}�_���/S��g����O����V<6��[�t��3����by��ùc�)E���f�t�&�u�1K�m�
������ �x�����g��aƮ���o^�X䖟*:��^�v����!Ҩ�PQ�i�d����Ӗ���`�^ ��k�z�!����e��4�R(k�g�L���X�$�8.MJD(}M�=�P@�!pB%7�/����B�p&��8���ٛ�^�-mKos&Gɨ�]�QUsͼ��Bc�[����v��m��Nb	s	�e���	�:��C��r�"������P߆
��	���MD�`G��r��1��Jh:��w�c6T��p�,t�a���N bY�� �2�p���"��[$�h�$f(�HXg�;Wh`��W|Q����qj�^w�����y�_�ؔ�Ȯ�:O%�"fn7. �v��v�	��/d%=�^{Z���ڷ��L�[|��R�[�r`Ҋ�~�E��Z��Q�K��)C�r(��2��S�����B&��J��buP��s|~�,)F�M�����t���#�nǂ2�c7�+�Y��'��'�t��:6_�Z���L��~�������V�q����+�d܉{���L��p�$���d���;���G�`9��:��c&gWO%ԼI�o��%�#)]C�#��U�Pb� J��E�ݝ��d�񝴝5��N�}��a�E�ˎ	�t�1�\8�@l�޸��6ƀ_TI�?9�_��9�H�[z�#��<��2�E�N��O+~q�-p8�]����[	�}K��*���f7e�D�=R|���Uڔ�g�v��k�o-s�U�P�FR�j"p"H�D����U��WT����s�J��_s$
�f�;���x0� q�S�6Jq]'a�e�F��z�҉�a��娨�G}�� ���5��[X�@���n �'�8澿m�,���]��tu}
��ò !$����=+������&|澡HY4��r��/���?5��o�TO�>�ݽm?����F?@k�V):G�����>?l�8��9�պK���C�P.��1��e7a�:�EyP�~�e���{��'�`�4焿bd��#��)�㳚D;��f%���S	@��|�#�Ȣ ���}IR��{�5iV�Y��)o0�7��M�UĘ�/�_�LT�/�1�N���;���}h���}7��+�6X��H�|( �b���)�@�S�˝��f�8�m���x
X�� ��1V�󥵁[��(��ع%��61��|�KF߃8��X�9���C��FRֵA��RMj�u�|WǍ4+̷����?R`�OieM�����nWsr�t(��8YEd���hJ�s� ��6N!���6��o�r�Q�;끹�d5���������Y�AϷ��,��2昴ҕ��s�������D/��`���͙�=���bx�:������~9;L�7tfǂ�.���|����0����L�D�?ʽ��s$��$`�a&��C�8v��b�<-|ÎdR�Fi��$�������
��	K6�k|� jq��q�K݌�Q�(��J�k����!MW�Lz'ҞH֞�#���3�����Qc�R��3?�3g�ŕ>�I{R�j�wc�-��Z(��MU�??�f��Ih`u5�4Nqg�77y��N�^t����X����r׹F}ј��F�%�.�v��XZ�\��q~ ��a��:(�/$����G����(t��%�븹�D��8�.oDQ�!c������]]���U�F<��h�c���eh=���		�n�˲Y3� P̊�=�����[�wT�	�e���.m�[��Y��`�hS�����ܩ��.S'U�5��W�Y����U����q�]A��l���TGO�Ҫ��wn�����
������7YF��wVA�_��bFh8U��Ah՞��ͥhq�+��Q�)i�Y��fy���r�u3B?H��k<f�G�	/p �@�\ ߽I�|��ċF��oQ���mY	�*���E~�b�������P4��#��4�R�*��W��F� �q�]}�28��L�-ZlQ��Ql�	癁�d��I_�=^0aj����\X���N�3S����P�Ɣ�y�wh�K��9�
��l���/?ӳ�t�~������&��i���T����WL����BO]�Ή3���	�+�tr��`�R+��i�0[M�
�$5�W��~-���no���I__�Z�iBt 21Z�}�ʸ��jc�#��".���҇�T���P��#���L�7�Q֞e�q����$�F��=�G:dQ��`됷��=��S�$�%��r�v�
,_Q�kgϔ�1pvI�<E8g��8W�>�P4ϣ��rl�}0��֞�{p*?\/�����J��Wޞ]&��W��b#���>cC� `4Ҟo��f����Q��%�	X5�?��,����S���g?�RP%��:�g�f J�g�n����	�1Zn�B���� ^^'8R���]5'�Q�k�v^��>h-�a��������>�GOGk ��,�<�-���a����WlHj����5�|N��>Szӓ7Pxl�]��Y[/��8U�կ�n���}F�=2�x�_&"��t>N�>�nK����N8��Ԁ��c��Wh2N h��r�חx�'
-�=Z��U���w$�#b��}�ݖ�s}q���2V
�tvt�.e����3 Y�q������+n�6Uܛk���ŷ��>��dN͏K�P}�0!j�W��~��|�2m���	��Y˪޻��
�;�le@x3�)*j�Ԓ�32���cv��Kڜ\�Wv��Q�q�kj�9�j�)�B�F#��@fۡMaf"�Jp�nh��
�������5%���c��̑�=rb.��vs�l�6J���K)GY[v��R8bAN�����CR�9ڡz��3^���?7�Br��a�?�Դr��:�\���"�n�}��.{z�_M�lqP���T�%	��N(��H�N<<Iv��E�B9c���5�_�,r��>�6��7���*�2�K��'�'{b�)9�L�&p�fY���}FY+����TVhQY�u;���x}n�{l��Իa���E��`/�HV	|�E��<w�s��6��8�����Ե'c�^�c��P�I��2&���# 	��R.>�w�4��qO���a��	��UUXc
4��Z~����U&UP�kB�g��	�$���r0��~9�e"m�Ǚ�E���`,m�\gho�;�<<���	��$����bw��fB^����ɡ����J��>p�|��N�L�(��4�~;�i H*��,d"�5@@�Ӹ�9��et��Hn�������_i'��Wٷ�\ddۣ����8R)-��ҩnϐ�岜��Ǟ�󳵻K-���G��������ӆB�3`2s��x3��h%�ؼ�r\K�j�����GǒI*����i�^7� ,�����-J�W�z}�V�L���\�l�}օ6��u a�;�UY9�ڄ ��hl2!�Wb�%U���}Y���w!;�|��ʡR@��5i�����IS�h
�]$��nr

d[����ƤrZ��H]�<��r����k?;���7Oe*���Q��
��	�4��؂�y���0 A{�q�}$Q���<�]a��� w�.Hmu��1"�/ s3�n ��ٯ�2���&��{4��	��L�]��>��
�bz�F���Z:��6�4ĒZ<��%u�ha��1�	sF���Y�+������1����A"���H����3��<������c�����6,\i��3�DT0����hJq����!�5sϲ9���I��� �G�b%�$0a�_�{�0��ױTo���8@��Y���N����M��,�9����q���\cjڰE*���6��j�;��G�������p�_jG�5������ؒ�A�o:^<z�-��� ���X�G�C��vCO�N�t�����`�?�������2�x�eu:���KI�L=8/=�xP�bM	�.`bS�KKS!C`����O����A��'��$�7�9��c�WHau�_��?�B3�k&}n��pj�_����7�Qw�-݆�pL�kqx���e�"��?xD��TNL'��4؟q��Y�����u��� �1��� =��8f�5�fO'��0�3�Xj�-}Z����Bh��_�m%��_A�iRM�4�`D�bs�~e�p��Y����=��剭��o��e��Z�KoX)�3r�)�֟�՚'V�D�h��(gW3-�7�{j�	���V�U��]`����$�˩��/�{VWJ5p1o�Q)uc��b��јQ�T�M�=�F�����ͭ�l�Y+d��H�8�/��E���ϝ��	����b.0`_� ������`>R�|Z���ه�a�G@���z�=����9�1� G.����9�Ӣa�?�W�����0�q0E�d<'mĝ�2	*��b��Ļ��"7?�7�vV�Q�t��jTm�� y�pP��Hp��Ɖ���4�i-&@,Ӥo8R���	�� �����Z5��.��x��_HtMo����G�"��3�hQf�@�1k�0�Bad�Mη�E��(���*V�Nّ�C6/�Ӟ���c�1R��s���LV6x\�0�*i�@N�H�@�N�/�nk��~WG-�}�K��k��xe�P�Ͷ����}�y��*.�'vN@+��v�{�5���˗co�,�P��{����#0���[G�����dEX�/WG�a8g;G�3�%\VoN��m�d�GW�Rp5��;bL,�e�o쳰��Ь�'��yoKm��ʳ8��Df0do����I#�g	Э���V&E��R�p���Q��|���̪��@<�sF}A]���,l���'���p�X�epia}�=7;_�?�LX�B�U7!6_D���������4�(�b`ΥR�1��P��r��BO���\��4�s��Ú�2�]�g%� m����>8����\�L��e^E�`uZ0�z�����ǚ��(y�N�V���w��ʫ��K欇Urk����	��"�Ɋ�9�e�>�d�����!:���w ZkN#�,�g��ס����9ܡk[m��Q����zЎj; ҹv�*Zz�~����w�)�I'[$��Vu�Gж�(�M��Y�A16@�������ӹ9�Oc�����`�����<����� ��݆��Ni2���j�QNdY&O/�s���n��K4#�$���E:�.C'K+�J��*�U�&�iIט*����a���EŃD����jd��
����Īz�A	�17W�խO9u���9�J�X����s����h=���;�ǁ��p�\缼)�ig�|o0#MQM3g�����p��6En��{�L��ڀ�3�����ò�m{8i�soW{��C��k�xC��]����iT��at�ev}���y4��*
g.��3�1�XMԑKQ�% ��Jk������W_9�v�W:��ۂ1|:<�~�D*7l�;�
�J+o��7A�Hj:���S{@)$���s���@�ʓ�X����OB��׿_n��{Ll"-�k��"�O<�ݎ�ۨW�q�&u��P���Gh=��k,����"f����z��F7��α�S(܏y�M	�mj��xD-�,�;�	�b,�D�`���M���6�+��[~�d(�q�Y��H��S�ն?]LT�^$��ɎtW�i��O�n������H_0w�]N�w�����wV����J�Q0��U�"Bb�xH���6o/�}��#z9"kA�'������
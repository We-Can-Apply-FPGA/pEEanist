��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�8Ӝ��'�����@OI>��.Q�w2�D�봊.������D��H/X�c�'���)c=R�h���ֿCC��,��5��>AR��#��;�u�G_�p�G��%����;0��N��ب�<A��ռ�c_�D�ȫq�-v>�?�'���5Ę�-�!��#��E[��v�V��D�=�Db_�L�>jGj��`7�+	��\�nL欳)1�E�_�h�5��9�U����}���n��E'/���R��^;��a ���t�'L&Bo��Dg,���q�vPb��{��/��9J�����μ�j4AȖy:��$h�g����(w�"Bԡ�W�~D�6����!�!Җnw��!���T�
3��niՓ��$dꔙi�:�F�}��&��Y�* �(�ـ�k�'Y�p�p�łY��d�w' ��1S��i�����/�߾�~�^�/���)`Aԑe�nl��f%�K:p3x�BiBs��+F�@k�n�������ۋ�X��I8#X���
9���(��b�]��w��Y���P*�����01��פ��B��3升�<}<���J�`�=��맖�ڝ��c���e���������F��'b�����dXB77�	�{�.y��������S0#l2Wʆ�SH�J�p��"�ν�?G��0:n9��� l+گρ��2� ~+���]A�lάc5ǥ�)�t�.����\p�o��OY;w3����65�������EL���X~8�/�r���
�kL)��FZ��kr�]'��J
��}�,f��#�=#�$X���A�b��������k��,�E�k{!�"�NS�Y�By�ř�r�2�4�i6x�c"Pys���r��P�# �^�Z���;,��$O��X"�[�^�z$>zQ���K��85QE�������(�l3/L5�V��Њ4X�R$Mi�l����%�Y3��2/�O�Q�o��9���d��6QFng�Fb���^T� ����-�	v�u��b��Kӷʾ�PR����{Q@ɭ_�a���ٺ[�m
�}?O
�xK��F��*�/��Φ}�<��K�M7tŠў�(�iȭ��M�� �~<�Oyz��sX%	c�>y�Nj�V0EƢ5O����Q0�����0o��/DۀU`ڰ�E IWK]����c��M����u�P��)�"NeZ
8��dhn*����i��-Oaּ��ݍ	p��D ��Uk��������߬��j+6������CE�D2O1�X=}��~ |�M$]v3%�I�� ��ͯ�y�]�b�`Sκ��Y%��� -��GتCHկ��
o��-�03����jBn�i�h
n���Q`%l<��E�Iy{��("�VN�}��A��b�ݖ;���b������������_����)a�H�L��_& S����O%���\�� ,�_J@ռ�Tp�DK�W_�K�&@;����j���X�_$sC
��n\b�mT,�X���@Mt,d�����'鹞6\�� �6��kZ�� ѭ��t���gP���~���"{g���{QL0���촗 �і��W�`ڰ�/GG���{ZEh�S5�C>T'�4�c�@G>�5���5�,��c��&�\��zR�نĺ��Z������U��A9�EV�.Bi^_nR�u�%ڐ��u}�	�㋆�#�:�*��F�ȟ�9��a�(�1>���y1F%Q`���u͍����f<��!E�!ܬ�&,#U����WN}o~[���7��c�� '���(OH�^��=� ��_J�+?���$�^���$Y-�� Y�C%���WG��B�����[�tC����]
�`OWD�g}$%�x�,5EfW%�ǰ�C���{�5)Y6�;�<�������7A k�1F��uN)�F�k�j���V���.�����̄�" yZ]⯚ѯ�/V���1>蓘��y(,gF^�����	|~D���/5j`�
�,] }�΄�0���U#�R�V�Tv��W�}��l���٫�2�`�?Uݍa���ؕ��'O�����d�h_�4kR�T�z��0گ{гŔ-�r���V"����P�����7w��7��F�)��Y̞�P��K �G6�nt0�FW�Hp>rնO-� U��ˁ?=��ڈ����jR�h�n/��L�?JmbQl�ВDauJ(B�_�x�׹�8��[u,�\ʡI��4TY����R,�6b.���~�w�$���D\A�i��Z��~����y���mLW"~i�W` �0�4U)����\{B�oO�u�6�� �f�3멠� �5^Ï�?���a��7�̮=��!N\ �SL�զZl.�T��6�r�{� ���"��sʽfh�4p�&)�i�0�`�atE)��!aK�Qfq�P5aǓtF�
2�p��'Cd��6�S�_u�j-��s�k��W� ^�}Cc)!;:�ŐEs�Ԕ\^��
�L�ACB#����I~C�ܫ���Q����f�K+���[�"鷒���a(,�:9#�x�b�E�* },ɴ~�RW�.�z]R�R�$�5Q�@�R�] �#	�du���
��]+vf�$T�pvZ�aG�Ø;`� �鵸��Ebp���FA[#q����rd��ۨ=Q�<nL���TJ �Mw��,E%|w��BS.�e�����^�0�����c�j�H�e6Q��/�G-��W���O�W�R��(s�#�e��vy+~�\;m{����t����x�D����H1c&H�h���^J@HP�N��6s����Δ�>#���!���*�Y=�(	�C�!���"ŋ�l~���Uu̴
<Kq����=�G���k���z���X¡�=d [�Š�J,���Q�> �i�׽e��Zj�UI}&X�n��}�Ɩ�E��-B:G����� ���O��tv�u�w'M���R2�֢���B��h�䬘��"%(7���Q�I���m���&���c��P����{���b@����*������θW�!g�A|�2�)��>�`����A8W)vPd���C`Z{Q*MM�Dڌ2�wtk�>	��M^�ݙ#�x:+(o��c#�h\��JbK`��H|:��a�2�������g�̩������O6�ݕ�ĔD�.&Lq3FQ|4�C�քCbSB�c�=(g�qR��3���Hha��L���;!j4�`�p~�)���@�l<͐ݤzl*n=��]	�[�� a� ���c[�`��i��X�����R�F���"l�e��oի�r�]�O�7�������9�KE��[�$�ڵ%ʺ��L��Mʶ� ��ңƎns젬sGo3e�������я+7��� ����^���_j�]&��y�m��	B8>�*ڤl�e���q�1��Z� @����g�+l���3���#bĄ/�+��0�b4RӰ��_LR��`�i�r'��˅�Q�3���m��m��\!&*S�$���_9qd����_{T�RH^�T�S.��}Y��JW��UP�!�+4�J�z~���'��\�L�"����̷2��et5#�,$8Jy����F�֒
/�V��cN�9��7�����XA+��p��5�_���`Tq��'ؠ� 
h�����PCj��UX�S��D�	L�@�NX�.h�{7o5]0)��=!�w��?�q�gH�,<�M��L�5y�IT��m�#o˃J��9�����ޜ�����?�	��,�d���?
����ܘ��fȫ��#��j�ۏ��é6�N�u,9�U���OXZ�u"(U�_W��@�k��$?D]�wZ����]�� M�#������f�%B�;ʮ.��f߬bi�]�*�_�4~�>�M?ѲԼ��6T��v�Z�'��O%�`���5��[�x�x�XW�<�I�T\<�F�Ͱ�[P"C��ʝ�}a��-�6�$V78���ANeSe2x�?�9(��������1NQͩ��]���r~tWVp@�ks���<�%M�,�mډ>#�hLyd����׾E
��w_�-����7-����s�l`�&��{��rk R ��)��b�#!�:��)��P��!ZX���k`��!J�4T��tQ����9�����S��2�A���-����ݚ?��V�U�|�۽��QSJ�l>��w�5;�m�ctl�_oJ�*��A��ZQ����Zz�K�#.p���L����w�ښ�1���F�R������qƀF�T���"cd�M6�;�)32�xg�MU6��Yz�o�{&�`(�B�Jt?�8�S�p�-��K�B(�4R�S�����A���x\^��+k���Ն%u�֓i��%�S��X#7�r=��ݑK�?IW���ynL������9�1s_�*�x^g�X�!�=�\ª{}�*ꛧ���_�����@z�����E��le���EK����b��q�[��y��%�s���)���Y�?��S��9�CuՓ��:�Ɍ�u�Z'��;�B�:�{���͈�FT��e�c(]ՙN�m_kH���{#4�M�W�6��]�bi�%��C8Mn̄�jc�ȫQM�)���لi�/['��� Z��(�"���mIL{Z�ߕ����#Z�MLô��,�<J�K
��4ٯ�����'54�Y���àg6�e B��~iϿ���%����g�XjX8��m��A�V�I���-A�7 ]�*0���nt���l#��G�eRF�o����d�	ß?A6j������QG�Е�� �1 �>]c�Q��K�%f�aP/`�O���\@��C��ƝZ��j��*�k�J��߫f(�K�gU����B6P��t{:��`)T>b���Z�_)�i�������<��7���̰L��
)����3�	�M=����q"��Th���A�@"`������;�`�)_]�����8��6���I�n�ïj]Ԣ���VL�0� {J�{�n��c$u.��"��eY�Sˌh��w�$Srºk��	��-;�a��|��̦�'�#��Tt�&������q�"�$R����u2����N����Ym#^<�A����x�}L!I7T�4ȵ1��?��Yݩ �琏��;��誻��xFk ���Ʃ���(9�YhY�e�)�6�%�#��hI�=��S�yB ��1��D���{"�'+�)~1�i���n�m�̥�0�I�0tvv�s��Iz��2O�����[}�8i�_
��E;��܄��iG}�
|M���T[���E�bѥ<0�uZ���o����i=�Fp��ȯe17�"q�^y����1�遮�xEh
�2ї2�0�;t�p/����\�6hHԠ���'��h�&F������ܜ��z���T/���~5[�� ��^�S�E�l5OF�t�9KnS���1rI;����5�ꯢ-i�S�0�jÌ�U��\5bw�	�����a�m����6��\~6���)Z���?��B�Mq�7j�X:�$���9[o�����O$����{:���Le���Ŏ���f��q0z�a�]�������z0�0�b$o�V{����rQ����~�$o�rǜ�R1.ю��&m���&�5q��f����r�Eϼ��ӗ��QT�i�Nb@t�NZ%��vg�e��X��Ƭ>,�]�W��l�-E4Ƹ��*���5��ͪ�m�&����ݞ���FTȸ��n-S��6�1N0|��soV�]�@ǼӍ����>.b��T��Y]����Qg�3�I��j��aD,S(r��7�%͸J���87�rȜY�Z3 1���L7�����������r+�W g�!El�� S���I��w^ƜЎ��Zc����	�� �C͊!��$	��Lt
���MH���	�ǟO��F�4���H���\�����&��)iK[݌[B����D���K����j�~�v$�K,��kS�vƺ�#� �!�s�uA�"�;b�/L9��Z�����v�KH�B4O.��N��Xw�Y�J߆f�(��q�ȭ���a�P9��0�:>�vj�J^���|�/��3�	""�/�P��h_�M ��R>��+@8�3���%ȐP'B���KC
#t2�J���&];:vE�o"T�����v��C+gf��)������`����%����~p�/�{�������7E�q^u([��W�V��Z����,J��l{���Xs[��CS��u��(L�.������d0^�����+=�*�}�E=z�����!��G�q{��MmjƮŴab�	n��y���by*�I����T�q�G|*T)^��4I��?�����������k�s#�m�+��7L���6�Eԁ~������`3aK�D8��ħ��o��+�f1pbV_L��m�i��l�F�xT2��	��?b�2���ȕ�/�=w��U�sO<}�p�������no�$T�3��zDq�ei֩���G�-�ؼ�@�����M���U��_�-/��������뒈*�k�ʜ6��*&���U��u PU�J�M.� g��"�H��'E�H3 m���;��eՓ�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��`Ղ���0<a6B��(I�izr��6����,��_��M�:��&�PH���da[��a���V��z��#��bV�#~Z�T�����K���]��v�Ÿ����e�Ǐ�U�F����XPd�}�4T���|�������~"�l�A�]^^R�2.���1ח��:bZ����Q�E/4:�He��"`�XM���xǑ�/��(^H��v6�j��2��F�爴���9�2��y��\�Ob�w��Ne`ӷSK�z�41B���٩d#�*����]�o�܇u1@bMJ�L��2��]u�:#�!̘��*|Q���24����k�)a+��upg�9"�bl@Α�z�y,���q4ꊙ��>5+��+�_��BE���g��:	�t��}3���T��o������)�4��szѭf��H�^����<gi�\�����e���!�b[˳	n�<bl�oDF��VZ0��~��E�!E��#߾�'!
�(�
��ڳ>�ʲ��;[�oΫ�H�cuױ������l���$�P\C\$=����Q�,;~���A(W�o� �$�Ё��xi�="�)G�:P>ui����a��X������&��[����cOMM�����=�X"�$�_#����OSQl�hP�A[�L�Ot'=H$B*j�&��+-0j�nV��
�e٦"yNM+0�e���ޮ�H0��=�/j�`uv��dF�^���D��w�D,ȫ�A��}�|h��xI��*���m_}�a�21����_������n�'�׹�	��4z��ʗ>���U(��5��`�W��)aRf;7lj�t���d�?4Z�m;�`��x� [���,��XnZ�rذ�	�O��/O����]w��H�+s;Kk�r�@MF0b+��3����w�E� ��ʐ�O�i��ua�����Pk���P��>�ա3�Rw<�W���\�5�N:�_���t��`,Ps,	_�a�����UE�7�쇤��3Ύ���>.�8U����Q���\�A��9���(r�3V��Nqc4��"�F�|k�І�v�s��-�)��Ұ�x��Rw'v� ��/x0�����j�Y��*>)�[�4�nq{`�H�:DU?]���M#�9{�0t�~^�T�W6�<9��vׄ��E	���P�n���b(��']Ǆ�h����:
��mI(U�T����=�:*2�8r�K���p1����n��"m�gj��2uJ���%NK�9!�m��e�c�_��۾��Tv9'~xmҲ�kIfE��E���)C0X�A������8����������{���3Q6u c.A����*;y��<��=�i�����x9#����:E��	�?������Z�щ4j	��H@�9A;A��=�Q���<s��ɩ�wI���%h�a/�)�󊃼R=s�ݔ"����K��M����s ���a_�&T���[A���������g��r���;��xIK2�~�au�R�*��Y��X/����:�V{#U�`{}:�9g`�����U��Ok���.���O&�5�� �-��(��l��qߜ{�ǋ��ZSj4;υ
u�$�Z[�!����G��EM������ٱ0�p����4��Vj��sKo��v�]�ܡ����tJ�=u��m�ψ62S�r��pj$X��U��)�絵^��탺���'ncNY.�`q�x?l��>�<ߠ,������H�� s����袞I/UTRz��p99����`��Ԝ�B´=�P�I�Z^OÝYs_}Hb���J�40�Z7��s�d���)jb�3�Y���?�3��y��'�
U��Rea;'0�-b�D�d��")<�RHv�.��X�V���	��f��$���C�5�2TU�N&5�r�U��@�������pC�uE�ߞ���F���2a;iG2ԣ�Z��e��ٽ���6=(��-X��c�w��QRy_�<t���q�$�O���M�ϙ��\X
ɕ�^��8���K|���w$��=�}�e*E�>|T�+)k��KvI��1р �
A����� 7V�K-��g�Xdgt�Ö�11P����P~^ij>Ҍ3��L��T���D��S)�@h�W�.��k��U9�D�h��>k�\��gvh��=���=⢛WZ��h��ڗ$���a��MQAe���]��ҡ�5m1� ��J��+��D�0�:U�K4>�L��\aJ����}�(W=��{|r�.~5ʾ���8r��Q���͔�~վ �Q�Td�2撺̠`%�^5��%�K��������|d�F���S ��$��f�Z=���FRI��#�%��I�.�̶d�[�U�RTyw�9cR/�p�&&��\����Hp��g�:X1'�?�$��L\�r�'@���c�]pN?+uI� ��B�/���7��L�
,�`��ݤ8ϑ,9'��M7�k-���te}_�s�i�(i�[�`�N>�s���_B�jN{4.��E��'t��Q���F�L�K��,ȕ��\�rITD_�u�O$}�}��}�rЏ�K�*�O�2DK���������?}�f�Y�J�f�a]:̲����3�AeYǉ�9,r�+m���j`7�����9{݉���%u�f��_|����[�� ��z-�B�cI���1��ޙo�P�/Or�ς���	���`أ�f釗��A �~-�

S��1ے�<GG��H%�4;���s �ڣ���P�}�.�j�zw`A���9!��v,/��pG��{t�1�DNǪP?ݕo������ N��oKS�S�����sp��+���}3������=΍�T�2_]�{1��-4��Vk��:;�A>�*��!+b��"�#��ڱD�t�	�G^nz�pJ0nR}^wCD��u������A�H���:�=�5���r�.ԫ],3)N׎w�a�A#��mC��r*�?s�e��B�h����R���U��}x�L-���6��7�č��k�uE��{�mZ�3p��2���>Wˡ���KY����H�ԗְ��.)1�����}
:ԩIn�#`�ۃ��e��y�7"{�C���s�28�~�hM����SOz^.bYT��C��\:J׮H��;�F��U��N8Z3(�m�J��X pyI}���=v�s���&�.;�҅����Z��u]�4v)f��h���C�P��F��:t�ȟc�1F�������w�+dY�,��NI۸ 5L�ȝp�%���r�O�x�q{�Ghڀ�D�`���B
ٖX`t{��E�LV[�&5����0EPWa��F�u5I�Fi��5w|8eQh��P*�ld��Li��-6��x��j�d^�GG2�Gt���y��֖�9<�n���%N�Sw5���;~U
lK\L� �L���@�I����P�W�1��5�+g�96�1�@s��������䉗h64���v�v�t4²��$�����M����]����Y��q����蕫L��*>�%T:t��?(J�tkeu��ƨ�p�"�xQL;���t��1ˎ^~��<vc!)�R����O���,��՛�`�i?́:T,���5\�e���8��g�~�7"�Ү=gx�P<D�����"���HW���,��z�3P�8!�u�Q/��^~�k;�8̓1eg�A ��F G��:+��DY�#���ViU�idb}��>�.K��ny��]�މ�ǂ%ĩ�G�{��8+��Y�&n����C/it�a�t�(�9u��~������f�i3Z�"7��h?���j��֞g8�5�i�ʋ �R'�}x�Y�B%���`Yy��OXH[c�w��I��z�r���,��F��՞$-i�5ƩS���I�I2�.�6a�ׂ	yH�;MK� "����(�t0�X��Z��m�u��lU�Yѷ��ɣf��0�=�]w(́R��Of�0^w�9Pz����c�r}����H�q�BG�{	�P���}�Pz���44�q����؄h��]4�)���I:�ɪ��Ie;�-#���ݢ?���&KHD�nl�}5��=��0��Î�Gʻɺo�Yf�0���ܪ]�p�z.�w#����؎�i֐���GN��5��!���>^9��Ζ��x��ZL:K�b��D7�(�x�r�����NF���܊�(w��}xc��M�ZQ����Y��\�0a��I;M3˚b�[��7�("L5,I��	�(N	��g�dK����p�fT[ָ յ"��N�m`Rb���h >n�Y����`�OA����駍����Y]�)`�?�-p\��A��){w�:��cH`���~�R�I��m�,CA.�R�2bz�}��a�q�$�x�"��?�bV/El͑����Z���PT� ���U����39\��(Hn�D9#8�&��7��~7]U��`�)rh���u'���E$���7�}���Iĵ�//�P�Ս�
y��&Q\�^�Mh��^(�%GL̺O��J؜M	��@�̏b�C]Oy��.��h���������}{*�i�R�m7X��w0z\��D%F,T��'\@�Zb
�J�j�dEE�H��p����t���.���p����p�#n�O��B�n5�c�}^�����fU�%��g��	���� {�5z\�ܼs�`J�Ix��f��q&K���h�y�! (F/9��Ϭ��F\F��x)�$$��H�	��^Y�F�b�x!��}�ǡ���������׾�\�e�t���c�X�<�]�W��#D�%�}�0�D^,��=����|��|ߵn�&�#�28�'�$���w�&'�Q[Z��6�+C��4P�_�P����\�)�ñh��?[u�42L�S����g�v�4 �=� �U�V�Ik�/]u�硵�����;i<Y�����XMm�E�=k}���abi^�<^9�͒Е���Z�\p����b$�q@]V��^3�,���;Q��n�(:�hVQ3��r,s+!ɤI8�+(V4�5����$������1Jȅ������C��BeO��x�4P����5� �"+�返D�L��C�&�W�̯�q�f��� �vw��qN�?8��j����*�z=MJp� <��
#�h�mû��#�����9�����٫Ŕ*s͇��K�Ϥ}9��"��Uj#ӊƣ*��h�X��c��'��K��E ���&�z�]3t9W�����_�k�*s;u��ߖ�pm��XaÒ�A}��?ud�ꡯ�neV�z�r��|��B��� ����N�z��F�޺E&g5XM=�,=�L�2�zTP����C�,��O�f�G����^X����S[��
�|1�L��~ǾX�
rG()��b��<�Ov �s�I&Ŕ����Se���/�M�<��7������t�NS�6RX���\yR1֯��'�(��m�I�v��	x�e����{�I�����%Okq�����zs��̘:�籼��M���' ��f2�E� S��&����K��$��e�@�q r���OJ���*�v%X'�*_bwG�mlU?�M��r/� `�m��&�4�)wA�1JȆ��ς�m`��ۼ;~����%�����2���2w�A�t�M��䤡���~Z�?b�r��-��w@�/#�N�!u����<��WE��1��z�t����S��72��u[���t=b����ێ|���*��1�c����Y�Py�=�j}�Tt�. ��M�VŹV��zeӢ��}���Ѐ�4��Y������6Zi/����n��Lj�	������А���D��t�n�Nʭ�h�q/1RgL&���b<=��AeJ��ޜ�HҲΌ\N1`O6ZL��i��t߆���%6Xыc	q�S'��*���x?���5bxv��j�8g�����.^�>8����7� �|f�|:�J
.�]8MD��R-��9��i-���D9�����,�dUqI~q������	�S����g
����r�l D��&�S�H���z����:�SI�	/������[� Bn�ya#�I�!gK81���9p3�6���_�0(�/=������p�S��> ����%k��.,�g
hO!��!b��!��d7x�O�0�A��N ބX�����������m�D	����_z�k�d#��e��WW`(��y |K_�1S���y��ݣ�h]���/��� �󜝬��C��p0nc��gZs6�\\� ��D�1|#�R{{#0"O�iӪ�;\
��=�i��Uc�!԰@�z,5���X8P�aҩiF��|�Շ���C��^	i��2\�ìV�Ƶ�������j����kY�>b��'8X�f&� ���I4YͩH�|�b�	��������7�!7�a�Hua���^���g�Jk�\�miͻ_x@����Bz����҂w�HYG�/���W-t�p�6+b���C�̅���f";�(c�5���)o-�6LC�W�T���Q��{l���zQ�R�\��,d_�~�;/2�*�D�C~��/�Y�5���-1ԫ��U؟(�jY���Z)�q�[��O��hM��aA�y�U0��a��v	�bs�F���@��8k+��X��C]��3�F�m�:�B~��%��ඐ-� ��s��wO�Ǥn�-��]�5?�7�熕��s!'k�8����"ya�P�ء�	�۬ǴŻ�LgQ����o�E���}�9��l����yn��7E:f�j8H�
�8�R�v�{{�[��E�Z*�O�����E�K|�.�Ě�i�p�Y6�]iy�0��Լaߗ��C��QHyx��k�R�۰y�u�;��*&��LAd0C��!�'$�܂�f����[��Mn�54CŲt��Ǘ.x�=�A���ḟG�w�+ߙ�n���6�����"u��R��2���ڠLA�J�"a'�_q��XE!�}�����`:�Xt�n<�T�p�	���gײrq�5�� ᮯ��%���f7��X��cC���"Q�;��[�o0a���B����[SY+Z^9j)Bsʃ�fӈd(�5(�ٝ��\�p��erE��{X�r6���\��n����1���xWfD�;<&��ے���oS�UL�U*=;�q �	�E����쾁��-����J�2��	�ͤ9�[�N��g>?$}Ɂ�!���Y3��=/�6��{ �JT�ҕ�YHxcd�Y����L�r�m(�PBnS���
!���n�ѭ?c����'���+#�h��8b��)�8�I`ź)�$]�/U��ݴ��`EtL�_�؇��͏��<��H�25q�Ͼ{j���&1�ļ^�S�ptl{D��1[bm�,�޷����+�FO������k��t��^�4a���,w��w���e7i(�X;AҞ��g�CP��;�;�M����0ʶ}���5�ҡ�e4aUQ_s�6��T@�=�B}�sZ!����V���X��[<H��� ~FAS���#�_MП�B�3&V:����J��K�#U/��G@�K�R��S�> �����L��g縈�5��������6��M�N��(ݾ1r�wvmܮhPY�GSQ�E��c�V�����e���4ҳ>��	k���N�|FO#�}�?Z���$��»�9��hBr\bd��:g@x��|�P"f�k�&<�e���΀�R�J��4
lhQOyC�KҐ�G�=ϛ���d`g��H���z�}�TÑ�s�?�ܒ��V���s1�-��E�g���d�
,k��|z�*)k���ڦ%�D�����æ�������6��-ð>y�aۑ�9���P<��TH��>�w�I�q��W !�|X��L�d�=U�w�����q��2�Bl,��9�M�H�U���U5�'B���&~i�y�2�����A����bT����݀O�s9r�>�1�����nt*i�ngC*B�y?��3R��E�9�wQӣr�]�?8��w���cu+I�����O�n�������`ֿ6�����5P����f��2{er�GeF�ht��WN��+��?�}������a�c�e�\۷��S�Df��L�\��ɉ�+�%�PL�x�ފ7�_
�K�<Is-D  |t\Er�h��K��xw��C�W����>T�m��̈�W���p}º�bFʟ�@������oĺ�g&IݟJS��u=C�����r��LRxD�ۍ4�o���nJqv��s��z��#�-�?ZN��09:�O�������@oH.�_�ٖ����\�p�Ϻ��"���{`p��E8M�3�CB��r���Ȥb^��cVA���J�<�N��_��3:��'�̗I�<�z�����[5��b�i�j@�-¬-~ă�Ev;Oq�F*e��?���'�Xv��*.�>Ҕ��y|4M\]S�#1�M'x�r3�h²E�K$!�o�qͤ0�� ��P:��|�H*|ZO=�@�־�i(l�y����o��QkQ0>�,�ʉ��#r�sԨ��!�K�8�n���`~Jw�BD�ys'�X����`�#��;	��KO�f��h���7��~sO�����S-|l.e���;ڽzLQ��>dwő�1���:����Z�/�|=	@�4��Q���>3�f�����o�OM@��R�W�k&�z�&�}2�>����t���e��>�7��H�oqm��H͵z����� ��3ּnț��(��7db� <�؇uR��؅P����f +4P[ԃt���S)�l-]q
>����WOM%RC�Ȱ����
~�N�/�P����lr�g�e�q�)�g�HS�]&Ӭ�P�r�#�օ�dS��>Z�E�_��!���;��!��#*�d1��Y�]G>��<�/�B���	?��ė?��L.׭!O��3�ϭ�l�#&�(�t#H_�����I�l���je�WG�jk���ʗ��!�a|�e�<���k�"���)J�U^�qC��Ρ,Z���~*#��Ø:��}2s��0n���ξ	?��p�1��e0��Ȝ�ipe����7O�u�h<��([��0b��\c��1��X�!1�_�J�77������]���.��Zմ�"���9v�;3���* �d�f�ޗ�����',ȕRp���"}�lFb�bk�a�vGo�����]ׁ	�<ʞ324�`g/m���Lo��Jgg;�h�
j�FwJ���<,Gz��X�fA�6�3�Yؿ�"շ'\��~s�oa\�7��ꃨ��p��.z�0y����'�1ЦB����7�/;�Q���Z-w�Z�)��Dh*�t��B�j.!�:�I�����U�a�YD�(+�8(����g!L���Ҥ��{J�߽�.�@��*�L���kE* �����Kк#�af%.���[�%�Z�f*�"n�x�w;`�4�J����*�G���Wkjhn2a�������16��o�5��=\�M�Vd4\ɖ��a����|��t����1�*m��$:ະK���������ʊ �Vh��;�Ե�L�G�"�G�X�Φ�~�j'�e_�n�Q��J�E|�5�Y0V���&���S㚷(��O�>�G������B���"'�}�j��gz4�ۡ�|���p;�D�?��J��.F$�)���x.�yƞx1И�H)&Xic�oea�_Q�
����pɇ� �.�y�7�x�k����k�3Km�W)������i�㯥F^�d��)��� X�k �����mq�<Rc����>�����vO᥽H�c\��C��i���%&g����.�ޙ�?C�����ZPѥci}��:!��G�	Z��%8?Jr`�B}��]��o!�j���(��~Yu�f���$�8ְ�\���P���7����J�e��VD�[���儩�����%���T��w�b
G������JR�����}]�/�a�<Wی��F��S}��\�M�f�@�^;�㍡����/D+�� &�Q}
Cn�zt�~o��m�)�QW���8����
�9.�8��~���x�v��0���5��2���T� �T6�C�Y���㗹9"U���H�v巯d���mfW��|I'&02��1����d5qnf{q�e�[��r��zv a���u��� �<�������K�|iv�k�7�3)��� ���`�/E�k�Lb�����#��f���=�`�T)q���R�^L�r1?��Q��k�X�9Q ,����c7�Iח����
���彞�,�jB���bMĉB���1�C��b߅ێ���Cbm-;�Y��!��?�O9���WQ�*7���z�N]��1_�����"���f=i$�-�w����h�^��A�3�u�ǹ�N-����FWE�~%X��s]d���"�P �j�>��%Uv��o����¬:|��U.�>�X7~��>�c�~'/r播�v8�~W�M�*i]u�Kfb��1I�ܩ�˭Ɓ��ա��ܮ�=�
�6ٕn �	����ߜ��;t"h�/� S�FV�y�W��ce6��GR��1�1�l}B0��SdF�Q�q����T����r�d9�"	6�z}0M�L��u�Z��H0b;����x�˯���D-�X]�[�ۗT��#i��v���n��׉��oq��Ў3��V��Z˪I1�5)�Tu�4\ffGW�p�ЕNgN�S�!Kr-�,�/��H2ߕ��������:�U��,��k������#�[�X_���wx.N�ν��͝F��ii�����v�i���V�gL�=�������%|�Xr��V�K&���Lo?M�Uy�r�E@�)Ŝn�u�4+n�c��~¸�q��g�Pk��� ]�o�>O<�!��u(,�p�٦[��&�{͖1�Z�%�r.�w8�c`�(��ڲ>��Q�����J��M�k�[��k0�������W�l��R:=n�Honv��
+ҳ=pD4��D�4íA<��1ZI	��`�z������m�&M�L��3����V���d�W���m���oW�9x]�S@(������::��冪��c�
h
�F��Dʬ�.I�#,�l�������C55�������X�!�8#���K�,��˙��W���5YY+"lN)c�``��;�����FC�?Dr�����5W�$�n)���d�X;��zL�X� b(�pe�'��X#����A9Aѭ�x��*���Zt��P��^U����O@R\vg��IV�#�֩n2���6rD�����$g �1������|c��g>�K��߁����5��U�w����`�;�q�D��E.��x�V�%��������h��7'���4j"���~��od���C֍��z���\�y҄��a�������3yt��2��]�]9$�SG��rU�Lq|o�!}5�굤2�RW��]��p������_�@��c�V�3Г	ؖ�f�r�&�MAB�m�$t��;��:5aq}�?!��N��w����)��4�<	� �����@�w�����Cb ������*{`jV1?��i�98���몺Hc��{���������H;B}���}���U�\Jr��_J�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n�����n':�l�,S>�^//��|�`j��A�ߋ�}��W�:�c���E�A^��C����^�3��p���a"R�V��y \�����߉S���7����$7u ���}.z����tHBrFKB���G!ţd� ?�S����5~�jތ�u��):����`±�x{��G����n�;�J��E{P�_~�g�BT�����S5rU�_+����ZQG�U��	fh�"�8߭/�����p����
�<�wE �ƞj��Op}t_���-�~7WIS�^I_ws��z�ܦ�g�S��9 ��@���"O�J��Ə��'��C�9P�"��hh�4{r�Zq`�8$}���=�;���ߺ-7V�q5Kݱ�g���o��oc�OW��)��k�u��t��RX��$�q�	>���P�4+m���q8���ޒ��+jD��K���B?b�	f���Q�]���=�D��d �UN�1��Z�ᗅz���D� �1��aLR.D�h{�:N �	�O������RY�06�o%�\\0�)Zz��)\���M���8%�ޱ)D��k����6�0��F�[�+��h���}�i�q�3�2V�țI@,��q�����t<��XC�4�5�H|� v�N���'w��������rǤ �MZ)�+6&�|�U�:B�M ��>ĝ�-�J
<��~��n�p������l1nV��V�ù��-t��^�V�	kt��6�͑���5����x�gi[!� �'�cY�x@��6t ��J�x�
�CsH�dW�`�ƫ���wR����6s�\H�a(L��qWt�[����1�\���$b�M���-�4��1�Kh��
�.&�V��)d�F���6{��u�K�B �Vc���_�K�[/��$��]�$޻c�X�^�Q��WT\X?-Q�Dr�f��1���ܾ�e��w�m�P㈅ �D1(ԟȠ3�g�A���uX�f�(�B=��lP뇽������M�� �wavxڋB�2W�Qa[Nz�b��~,<�@�QP�A�3%�: ⸹Hð�{���U(�u��;�lї6�#q���bԯ����-wc��ȑG�s���S�U{�DvA�~2���ϫNQ&˲��a�zMz:a@%�Nx�}MHt_�*�<=~bܬ��m�+�jzu�|�g��0xB�������2�c�.��>9�%�3�m:��x�����7���BrmMńPO��ߋ����v>�V��@� !�e�z�I�g�UH�"��j��X����;�_N�i�^�J�����D@��C+ctG���f~���B����wF���:	���3}������
g��" ��
��#Oh��=S�	��P�e"=^�#m��l����Df1�G�u��z!���Blr9�\N�lw��֤/̑���X��Ag��ת*I`s�wT �
��?<�ߌ������4��|ϙ��Μ)�|��$ީ��T[-U	}��6�zQz�$xJ��-J8<�W�rـ{���|�%��i�CY o�T X��q��6��a(n��֍��.�{��P�7��q�O,�rK��1�vt[RN^��?N��Q�8]3��]x�5S��O�Oy,����J�,��w94���I{*Lڦ�����Tql�>�#y��̩�c�2�{D�N!1L-*`̙�-���(-X>��O��t����4���w��Q������m��оԽ��U(S|��H-��b��+}+A��%LV;,���A2�\E�w<h��5Rх%x����q��^�1�6�/�7��|PTQ/�?�Cw掕��*$Uߘ�e��s/�
tZ �w���wkЫ�Q���9�p� =@|ʞ���i�ĸ�t��:���.�Qq�8�ȓK��hB��f�X�ßj�m�G緧tQ%�W/�m�_\gs�3
����a���N.�'�a�{aFnW���������1an]�65`��
��u��!���:53�zꧢ�Uw����9��w��|�;rɵU?q�>$f�Fv��?��9`Ms���@ڜ�.�
r}P)�(@V��s��n=����6�c��,��׹&u��K]U�9=�d'�9^�RJ��FA�J<�y�c��CiP��WiF�L��r2�V�¢q3:�Do�@D��k2�\�����>R�#�H ��� 6z��aR�XOs��ET[�x����$��`�7��:r��If�'te��WR9�?##��U���o{w1F'd9�(%�l�PԷ��j^��B-��X�k~����Z�r���C5AT�8�HOn�X�r���)�K=� _�Lղ%_�[lМ�oP��$r�jl�@�!�Zytyz�9��6��,�L	���ʽ��k	�,�	�:9ķ�wU�����,��Β����� �j�����&�X.q��Lc����<�c��J͐���_<��n҉�ď-�h��IJ��MQ\��r�_p��������L4�������ߕ�޲���b�d��$I:��_S��q�Jyo�5�#��#�CX���$z+XN�Y�h�a�U*�ʅ��iU.#(��-�SS n���baI�]p�_/	�1k�iG�5r]��x�@8$&(��I��m;�d��܍|v�{>ef���?~�G'��9;EHOY���u�di�L�X��������=�܇aq�y�g-q��#�:A_f�q;����	ȭ(L����щ����D�ڏ���:_=t�͒��S���0U�*�=bS��>��!tL��+Ut���cE1)|꠽Z�uS5�,�[�N�jA2���ϛR@�n	�Y+l�!�y�d �m�+� ^����c 1���0��oێ�q�����a��C1���q�}S�P���w�I!��>C8?C"O�۬m`	�j�h����ԝ����82L�y@�'f��"���=��2�:��%��X�J.5@�rvz�c���`��G�
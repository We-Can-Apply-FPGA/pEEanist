��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n���QH����Y܎fy��no����4��
��q��X�`����[Oiw�ɖ�pTO�X~�jkݰj����TZ��� �m��v�s�	�wpM Ƿ�^���bxM�T����;��ý>D,R�XR�9�G��e����9#�����?�ZB��S}�%��;��ñg3��k��o�z��9E��}��<�Mm��t��.�KL��6d�
�j8�Fw#���{R��Q��|���J�����iP��BB��Tj�X���N��F��´��
q�"~�| -�흒����`��H�;�r�H9����.~�JjX�.�������R4 ��"�D^�k�fr�7���k�Rު�p��,/m��b�m��2�G�6�fe���I�%^ޯ����,;A�mFə��o3A��%�U�pI���Υwކse�d����%��u>�����Y��j�*��J1���v��[�iX��\�W�Y��=֡i鍭8��s����<#���0��Ѣ��|
��2ް�G�� ���'������
�q_�GGI���s�	n\��Uɬgil��w2֓��2L�� ���3*�:ތV�����ۡB�/�JD'߇�?ӈL_�9{�78!{cg2Ap��zgG��(���	�`���$y-Y}*4�b��E\]���\�i�g��
�l�Ȱn���%dh����vB5�&�&�G�~S���~�`�D���H�Iɱ���\��R�q
IU�!<r�c� �e5�E?�=�[{�A�5(�1vY)H����Ȩ.�*�������'6����:�C��'6�����_�����<&�1���!�5���v�+MZ�&�4����aS��.uxGB7�͋�
��nBh�_�^���Z�)y�G�f�����åT�/0��<=x�H���i�؀M��_-e��f]`���0�g�*A��Նs���H�Ȧ��1�=��ܗ��AO���7SyM�+�w�7y_��9t{�":��q���
�ᵚ�ih=�|�&��b���~��5�-5#��-�2rBѹb>�+�6 ���H\pإY�PB#ͯ!��XO5D���)�祀j(����ג�A�lSʏ_�������O]�"�^�M�� ���.u]�A�SE%,=GwE��E�d;��
gŢ����d�����~�bľ�bp�����2�8��X'�f�ws�r��=��%|�g���%��E1y�Tl5�ƄqETb
|���-�\��!�Y M�/���(E+d&CV������R�z��D^�e�#3Cr&��M»Ks��ptE��X�>̟Y���r�\��@bP�	X�vY/W㑒o�?�qؘ�x��;k������>��ĢS��(���	�=�Ɨt���.��3u�cE7��^\/P��2 {��"j�ʂ����!��kH�K��R'��>>
P$���с�i`z�s�Gl���UQ}/�a=��a�lpR6Tj�4:2�O3�$��o�C���GD�n���Q['�����U;�1�9��P},{=J2m���n��ÅZW�>@�*���y�CU��=��Y?k�Q��W�`�7�6�!��8�
��V*��$���+��ׁ�po��w��l06H]/�t��'b�����L����Éh��cn�/��z�?��W	_C�z՟&�7�c�"�>9�tz�C'���+�� b�?��3h'P��'	^H:�_�
�$���e�"�3b�1�����A֊&WG����Ɋ!>�\�Y
&�'ƒ@.��l?^�xk��A-�緌��ա�P�\�K*�%�ǖ�Aș�F�>���ge�v�%胫�;�����cX8B�	�@CQ����Cҥ��f��#;h
�Gk9d)�������1Q0�׉.Xr:�\�g��6[r�y�%�Њ�� n8��*鈟�<G��q��g��׷h�%%sE�ќr[�y�a�J��jw��J�BwBɬ� �}m� q��Dh�s����Q���P4,��H*��{?����)}��n��߁U��^D�u�J2�O�~�ۋ%��Y��sR����C��ԖEƅ��W�Ue�-�b!��.�j�� V=�6���S����8���0̺��"�#\����^� �H�����N#;�|��?����RL��[�~�e:������>cI�}�n�V1�m�Ŏ�ɂ�F�r�*�\�fn�RW��/�3	D��5��ftY
�4&?�OG����T�V��N���h�O�6�$f ��A��M8䨷�2�mU���]�+���$�~Ju9\P۵���~�@0����U��]��9�a�y⻒��w�h���92�T�����!;����#�t5��
��}T���g�� ��a�j���.�Z�\?M��*�k���Ҡ٭���x*R�|����8�n檶����r��Tfw1�,r'c�?9"�i�q &]R+>�i�Jߐ�����Wy��e�NQ�>e`���}�t5^ϧ �UM�U_�K�4�Ŗ})3(.fXMʫ	<M��'c���@Y�ܷq毱vk�hKH.����2��i5p:���X��<CJ�G�+sb��UZ6=��}v�Dq$�;�3��Gǡ��(i���k�i�f���=t�u����%^lx�s��:3�e�.1��K�| :��j8ꕹtՎ�qe�}�����-�K�T�P�(t5���^6	����Ja�H��S����_��d"��tyٰb���~U��_�5�/u��D��~���W|=�=�7�@,�[}&�
��1X>m����Ġu�f���+z�й�׭�ŋ(i@�ǣ
2 �����!3������]O>���:��jyi3{໌#DR�3�JnBQ{r��y5,��8��4����`��MAW��	%�ڛ�_z�UOSz'US�q+G�����'�>O��^n�C���!�c���QoENe���P��z�n�.������`;��\�3���΁�>���U�Ou���(�&
�Omْ<ބ��>����p�[�#̕����%�z�Y�_���v`�q����b �	Y�8����6!���-��5񾌩b&�Ӫu4�����C��7��r6����d�A9�g<W�=��}��mu��ўhGVL#��������&r�h!<�f�����ߘ�q��v��qA��oD����T��O+;���+�W�B�����8O�c���&?�A=��H�&�E���pP��E=��r��7��݁�ǒ�A��r�k�r����x�����'���6TKHUu�6������(b�="��Ց9A�0�c�������ŀ�	m�(z�d�p�?����"��1?�y��\��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n=���U6eI�L/WM72���"��(޾A#\�ⅽ�������l��t)p/�hq*��Uâ����WB��q� h�n(��>�G��T�Fm۫N�M�x��{iã�Gr�7Yg��D��x�E�1|ͩY��hȩ�h�i�h���
_FL}�9//W:�r¥p���F ��x�����O߹� �4���.��{��w�Ć�-g�MA0�犮j�<��A� 9�(0�����)G�3��6�
?@���eɻ��*�QX�;$sy��)B�Oy�#϶8�c�-T�J�k[<K.�Q>�����Ud�C�B����o^"H��٫���5i�D��}7�{*��L)_=��v�pz���,O*S�s]����<�u.(�
7!�9�1�/A�""�<S:z�}��$!Y;D�;�0�uO�� Ԭ��b�Tm�XMig��UA~|�(��P����yWc�l�y�����R�M�B)��03)Ӏe��P�7V{��3g���ŵ{�<a�}�r�L�nYiv�a��#������O/��I��Q�)����u�DM�,9.Ԩ����ϛu5�L�G=��|�����of!��F}�إ��"���J[0t�/����r��８��`�
��7��_��}��`l����h��d��z'{N3$EeWo�ui#���¡N#O�T��sI�Wp_o�_�˒����MWdbL�S�1h���6;��X�J�C��)�BC|ڄo_Ь5MKqDAr��|kW���3~3F��Aqe��AJߍ���^����j����G�$��t�1�"]�6�R,�k�Ǹ�<���MW��8��������m���Rv�"��c98��5�1%3�~I�~z���i4�<6����(⡗4'R��9�#w4��[m�Iѭ��D�`Z-��{~�Ou3��[0(i'e�1��tC�u��>X��tc�6w���F��5cOӠ;>��fj ��K��X���dꎇ� :X�[p��t[�3�ͦ�W'$�㘎G�}2 y�Ѳ��Q�����[�Y�����kT(�s�l��������3�]������ ���gm����>D��? ��
lᦽGr���pފ����/� m^�eN��*.:���) ��_��D�΅�6m3;�N��`,��3��y�O�>�]�a���ۭ�E�݌f�5��v��c[��J��ݎ��gr_�h)���1($fiA��#Γ+�=�9�`)E74��KI"��Hc_-�P�z %(�#Gb�\��[RW����ԧ�鴻�L�K���=5����s���:�>!0o��m�?y�:�-��mvצb��G�E��`������R_�]�lZA�(c��x�Xrݿ�@�tT��8@k�}���5���:U^m�lv6��y�'����މ�ڡ����Y:0��/;��Vl�#b��=��Z�,$�a��\}]��B��YЧ?�>@Q��1�9>P��S=l"�k'�jM��SsQ3U�lU�8��)X�爱y�x�]�n)�/�&�O+���T��
v�+�9�8ʂŇ5���ʔ��T��Y���������z|.n^ ��@Ƥ�:^òo�1�A�7Tmv����T%˚�����x�7���5GJ�V �=�:�������C�y��L���#�=�A�Uߢ��*�a���N]d�Rxט���oOv��q(����C�HȄ8ގ�X_<#[���R���*�ƙ�%f�F�#C�":�{���]G�ȞO�D��b����<}CR��y��m��o������I�FL�	�Ѻ�����7��3���FU�f����u����.Yդ�@���{�_#ݠ���1���76א)������X��-L�MDz��}Ie��w� �a�1�HM<]^�W�~��b���凷W�]J�<%_�0w7I�&�R�!�����X�N����R����{�?�B����*2!e�+���+|��d�ĩ�\-e�z�w�lL�2f˱ٯ D�`���"��e��]ܧ�i���w���	EqӮ:�Ђ4��$'*?�G��yI��#���XHD�`%s0� �S�����_bd���*qAظ gWo�bA<��xߌ�/�Go�Y�*����ӣ�I��C0�`V=ry��TA������1j�e���跹�~W�)nb����R�Ag�F|�{�Au#h���\�H�2�<p�Gem�Dm� {P��/��7
����0��q�z�F�_y���g��Oآ��gJ�R���lO����!q��M��ӏ�\ )�3uߒ,��j��B^3v�Ґ����t7
��0N-��%d&Y�`Ł�9��h{�)}�b�Ŭ&#�70tB���B���
D���xAm�x���G��m8�o.Qi��S,��Feg%n���%O����T0�����p�H��fj�y�U�q���h�9G�]��ug�ڿ&/h�;9VOR���Ϡ�g�����3����|������UaՆ�Iy��L�K��?�uw$V���2�Q�ٮx��^_��AU |D�Ss��������������N�I��L��f\F�$�iEfڢH�T�t}����%I�Fto%��������J�+���:0�T��Uwܯ�d|	}��S.W�� �g\x"�J�̋��¦���u���A{块N��;{&�?�r!���2�0�B�2��_d"E��`��4s�uJ�j����s+�:�w��Շ�C�
ף�v�(,������8!5�R1S9�-�F�U/�%� fe�3ޡ�ck�SvqR!a|)�&�!�T堣�-���X��[��Ҋ��[�@4b�F�s,�r0�gʽYS��$��pW�(�!�O����_��^��w�T9����B_<��p%�����H�݌B�[%��Ę�'<��Q4���:[ ���]�R��
�Z"]�o>�����9�p�����$�o	��rzߟ�㺧���㆙}����S&D��>��T��U�Y(r��uD{Ⲟ�j��_j��h��[P'l{p�w�
h�2`3�Z�� �����`����G51An�X]����g_B���ff�ՁO��^d76g���?�Q���7�	���*�t�xX7}k��l�d�@�M���$RoR�D\2��IR����a�����LõK�ER��y-�����R�r���=�TsǮ���pن2a�>�S s���"���-����P`��M�F��_� g�`��{�)�Z���k�ܙHB��Z+�d
�l�h<4��㩄�e l'�9���mU��zr�'2 ��~�t�w�is�����BعM���
�Þ�%w!�JLi���ՕY�n/Gi����	�^R�(,�bL q3��0�8���r3�2�8�b��o��>L��Q1X3��B	b5W�!��MU�V�4D@7�hLފ,�ܶ�GD g e(�X�͙��[Π,�ܝ_��4hM���8�?��%��6ɤm���'|?GGwD�V ����)���YXg��ljql���Y�*�v�N�\n}\�؀�M,+*TɁ�(S�5�W�j;T_�����Rm��5�'�k����(����-�( N�_�9�b��>�J<5��I.��X�q��Ǽ��]ur���dUU�|p�n�]uaf���8YOq�K�h{?]��u��߀
d����������PoEJ�<9����b_=�}�z�,O,pUHC���b';(a�&FXZUA��b��k�����.��'�69۶v�?sO�6�F�2�$3K��Lх�d�y����$�hP��2s� ��E�G͆~�Q�G�um�/��1s�S0���Bd�K����qƪ}h�_t"F�t��l.�,�<��ׁ��W����Β�R��>B�����ך�O�H���׾���~�-�EO����.C�C�Z�����/���6�#anL+�'y���)T=ƑT�@�>e��WBt��^�%Uz���=�$���Vk��B�<�An�n#AQ�JF#��ȡ��d�����MJ���ssu��,����%�Q_��_�.,d��@
褙�Y�rN�8շ����>n����*�X�4�>!��4:�_XiC���B�~Ć�mʕ��,W���Z<�#�<Ï��K��xg;8rkV��j���0ľ'b����ձA�c��]�鞾O,�w���^ U�9�m#?C�m�<�t�ANE�#��Y�z@�3�O!��¥�r��3/�L�Q�"yc�����9'_�K6��[�!��ԟ���E�+��(��)�m*���N~���m�x�#	C�So�FDk
���s.����2	��h�d
���a�+:�fE�j<ÝzN#5�04���vd��/s'�d��;Vh�`�zN���:�%���e�Eш5�P�̾g�� ��d`���!���U��������Z��.�2�ϳ	��})y��1�=�,�t�W��{�Vp��s�mV�#RKF��?�>�%N��p��|�>� C�]�Q����=�a��������E�%��g7vs�i2� R$�)ӛ���ʹ\Sq�j�ϳPү@>aw��_x���]��V��w�2'I�3|[�vO}<FL9�������ӎˤ[�q�եE\�.�H4�����?�m{��}fg��&5Yv� �o��@etqX��(</�B����$�����Gd_6X@x�Kd��ۓv<&��b����X�9�2x���*��u��־�`&��c�"v=�{�d�����Sܵ��qxƾ��!��o)tc�oF��|p�NB^�	�%� ������>�:�C�����Ǩ3e��gdU�tp�={��Sse�H�w�B�X�Ai�<����~XE:�;Ld�Y�htj�5���3�^Øb���g�4��z�@�Z8����?�%�(t)&�(R����؃[�Ԛ ��w���;C@����Д)�F#��Nz�F�K0�\���L1���hŎ�(Zk)�iQg3W(����5�c���{��wgU��E��p��j�{:{V�x6�̾\�e�j������>��.}ֶ���ؓA�vr���h�O�ݤ�\3�#�Ff�ލ���8�%L�,']Q̓VQ�8���6Q��`�ޝ�Є������89if��L��W�vW��āD��_EpQ�L�Ά���{�a�O�گ3��+Pp>]0��X�ޗm�Br|Jc*�@]���l�=�x!K��1�U���b��<�r��>�ҽj1(K{ޘɺ�91#Ŧ�t������m��	����b�͠��}Igc�P�`���\�E�0Y\
�z�T'��2 �<��gӴu`^q���H���Z�#�6���i���dsn�]�W�;�¦Vdd�[�>LVÌ/���t��S�3z�c��<#�LH&�_�X���Y����ZE~�l���a�#��Q��xD�����q�<I�I,$Fn.� �[��2E}��x�1W��a�l����F��� �<�W9�=�C�v���7���uOls�mВ�*Q�g߽�A�rUy=�E�K����=L�:B�*�(�7�Η������#|�kE[���'��f��/�F�-�������l��zkg����O���
��f�g��5�yq���o����)�:-��.��p�U"�f/��K#[(z�
}�]�-]Q�Œ��>�FK�rR�C6G#k)��d+�k����tF�'Oϋ��0t��ԣ+�l<����{���Fŝ��t׊�4,-Ā��e'w ���+��6D�bʗ3i�7Dz>k��pҿ��j#�
*��	�"2���z�:�.Jӳ +|a�4�~��WO|��E�Ά�!��x�lS��CrH`|Z
[f%���w�b9�UFa}yȳ�j;���rx����Xc����tlK6R�2�F����\��඙��N�W+�Nvl���y_
�\�P�aE�;\��Z(��$��N�ܜ}�8�Jʧ�����ᣀӀ?��d�ӅY�GK,w����LV�{���d9ON}ս�(p�픦מ�Q;�<Y*���N����hjX��<MN`��X��|Vt/&1��o�^gW�e�5��$-l�(z@�-���y
fQT�_�I�F]�27�c8.� wivT �>b�PG)%6�� '�C��v�[<P1�xw�Y�����iM[8oPD��]�4M�&_.O����qL�D���1�RG7�����ft���OjV��{��X�D �铿[���d:Kҿ_V�jv���K��k(+9��7�4.�Z��Hs�u0-��~M�	�e�K�ËJ9F�K�֠�����B96Ga9�ȯ*j�"3���	�*v�fI�V��cJ��k7�(^���X��I*�Q��q^�tۧA���.�ÈH����~ߓ�w�����ֺߚIχuNk�0�ҊP��sA��iZ�BiI����*��m� ����sB��_�,<
~�b�̑�9T�.�;��5%���\�_)r����"~9��O�ioh��oī��}�|{���`=�z�~�,o�R��ӏ�N�F�p@C����X��aZ�=~$y3j��?�@�r����6��S�-�,�p��Lu!�:ic�[R<v�0���Fh����*�;RA�"p9+���7EXe��bx~��	�����n0b���N`���oo���=X����)U�W�2F��9f�f��T2�č�2C�ϼ�c�vng'����9vl���p��puu��3�z�!��T�)z�9ܾjl�Z�!��m���@Ӝ�SB8<�����d=h��m��H]��"�ϫS(������ŋ#�OMn�O��|,�`�+$t�Dā�j��A�X��iWuecAG9����?iQ������I��|��̱��bd<��;_{��u��D��x&Y�zĹ�)�:��y�,Ϭћ��%�M�4��L�7�&�I��m~��}-�Z��@-چ��ǉBz|�v�pG�� ��8���<#�$��K&���3�����Z\��T�:k�{<W�� �8���mpDX�Q�=uW���������i�e U
7v�VV��e�!(fG��y�	�_!2�5��-3b>E��>9+�Wf�֖S����HZ+��S��4�x��1ąaa}C�I�����bd���9� EL:b�t|&I��I�*�S�K�z��ў��w��`�] �f�cɿ\��0��Y���U�z�xu����k��1M���Q��%Ԯ�������{�q��O��bl�{;��β;n)�qB�15��+@G�;����;'�����9�k��vn�����l��y5S�L�>���w9�5����2bb����A�3���O�<�Wdv�"�o�b�FaOF�F�z�xU�����������z	;EV���(:�ʩ3��6<��p�$c�N� �
�g��cH�	O-Z��2����\����X�����=c�]�[b~^I��:2�A�@t����nb8�&#k�gN�U]&JX���i���|���~5��ȷ����/p��6�S^'���$�D��P.�(�;���hY<�匐Z����b�jyo����7�Cb�W�����s>K|���f=�>��Rr�z�dQ����\�(�� O��l����D�[h}�fHA\�CD
s[����_!J�~���t�$uX5�͚�e*�m,� )�eҡ�~ж�]H�7�V�\��'�7BmJ�������|�/��02o�X�=����M�`�zDIT-}��SK��F�C'������qՏ���2P��tBwӨXP�u��H2��F���_<�o֯yW�ą���R�Y�nzZ��um���o���,���9��?�iw�<��������O���e��n��A�Q�^��k)�?��ô������vi g�P@��N��=��?����J����r{G�R�^k�6�=�(S2a�dڀ��=��B�LM��%�c?�#^R�l�/xV�HR?��Fp�,L�E�SUǟ����VD�b_㡾Lw[:'���6)�#���%R���wD��8r�5_n���Yx��7f�DNĐR�OS�kc,�Jb�=l(9�N��C�E�͇����{��C�,Ϊ�.� �Y���jx��fP�=� ;����<���
�W��2@R<;{Gz��y�_�%p��V4�=�K�{�7��T#G����� X�c3�)X7vJ��jѽ�%��{5TLw�o=���{�/�C��QA�X����S�ՠZ��rt?�Ν�/��Z�jp1�k���'ME�)��>M��^���>�4�u!�r�|$����3W�Vi��/+�t�,#��>��X�B�©P8�m��&W��U�7Y���\˥����=A����)Q�G4_Y�'TD/}�uDB�F\&�!���:t��_��B��M��gbӭ���9
"���o_Z=�����#Qia�_Q�\KWͪ����^@�tYZ�~F���Y2����u$y��Ī.*������}QF6�1\xsǶ�v�{��Ep3_�v�n�Jm4���ׄD*�G��|�t���d!�m9�_H|��oT�C0�Y��T��9�
��� ۚ�Ï@idϬ� ^�n�+2t�Wȟ7�t��]eI��;��zN3�`^��$qN�HU/l�tQ�n� �y\N��j������'QK��J���[��w���h�`��a������kH����[��ƜO���ĸ^�k��*��03f&���� @W,hgd��s}d��j������7M�&T]()�5$^�7X���H,x��}�#�|�0jp\�8XH��{Lm>�*�Xߊ4�`-G��j�A�+�Uķ�%*:f�7�$� �� �����+hB� ��JkI��q��Z�^I�&��Tu�h60�m��G�~?�a_Kw�ЖsFz �_����)����m1q�������YY���?�iU3;�<��|L�RG5�+5!pKz�J��U�z	-*�����A��-_�'��#V�G���KCUِa8I�^�˿�S0yd��M�� ��Bb8�E��=�&�;\��-:u�fp\'�����[ւ��7C P�!ډJ���#��^-XߣF���Z�G&pF��,�ѝ���L�*R�Eww�X�ɹKh^�E�3��j�İX�}��0�o�s��eN���~���18.�z{���7ϯhx��
��h#?�����t^/�s**���%T �h�X4,t�ۭu�Q��S�����y�tں���b0)�Y���&H5����ׁ�%Fc�����k�B�zp
i���O^ç��P��ƾ�;�.��/F���u:ç�G�c�yH�o�|����D��+n�:M	�?S��z2�� �˵Do������*�&)b���c��A��ċx�lfzC��&�?��uS�V��[-JfK٧�VƉ��Xְ�t��X �`��G���DP����G�v<��a�L�k)�[��\rB�7z}������
�������Q����[�����vڒ�Ʀ�X"�(7,!^?��W��k��J��}m�����U9���}�P���ݛ�}��y;���ANGo6 �㼣�xH�0}�_+Lhɇ:���1}�yI�^F�b���t�a�z���kV�'
�Sd�E��X!��Ki�~.�5-`�{/Ǉ�7�?Q���9��6�d�1���
k���b���Z�Z���.��9Х��1{��/��b�N�+�o��R������W���D�~�7I`#ڝ8/�p�������2�	X '*y� gҼ��f���a��KK�ʬ���f&x?c��I���:�&�~N@�n��<���X�������c���օf\�%���}[��wUg�""�|���.�,�6�h�Z0�P1��<g�|d�\jATS�����C��\�E�z�fc�s�����]α���R���U\vô*�kv�\A6��ҡ�)m�'��GEE|tؤ���� J!�UOdSJEr��,f�zg����k�b�0&�砮�!�n�����8^/]�˖�.H]�o�� n����c��Fh���g
���O����?���9�z����&��Y���79�i��>�M�h?:^���a1�hRs{Y�R���B�$���&Գ�ɒ
��{�}�ji9=�XT�y��&����u����UƊ�4gq�[J'���"%��ܐ��6{�%}�����y��A���˃��gV���W#�i�9��-�'T������$���n���R�1-}D�r��Hh�-�K1�Y��S����� ���{ࣳ�Ǒp�j��[VK>�G�rS"I����~�L��21��g�^m�Rd��ا�B��uw��4�	����E�۽柔3��ͣBWћ.B�痖>�@����D��LF���oL������9���ѐ���BS	�J*5S�|��O=aO�ۚۚ�x(!����q�B�1z��r��5=�?�z`,#�r�0�ɀ��tX͟�r���v�%]f�z��Y�������A��Ȁ$�s8�׮u�m�E2G�J�1�4n�8�{������ٵÒZ�W8쳈��x� �D1����m~!�]�3�i�[���=������T�1;RO�u�����-�������B̜�p*'c�!iO�=�	6M�����BY`�J�'q˹�����j���C�;�����h#v�Yz_��Sj۫���V�y���1m���'R�YL�AJ#���R��[%�ߋy�$�iYʋ�75\1�Ab�3z�|g %�Q��y�QQ��u�\��9"&:䆆Yv�&���T��v��-[���_�}o� i��3W���,�|b
�s��C�K2��A�?�:|����u_޳;н��&0�s�#S*h-�Y�-�w^xo5E��S@���ZrG�ٹIN�=}�4�i"(FNٻ���%�F��e[�P�
��4��(����G�.��G˘%CA3�8[���h�x�+ֺ�*��`p��`K��AyǙ�]�QF�I2*���O�O���Oӥ8�1�� ��[~�必����
g)Xi�l��<�Ӳ�e*a�˞7�Ǟ�}��Sr�+��N����o�;k뤁���B=��tw7��0$�WG�
�ER���G�+�z��!�9�����(w��n�=�P��Q�P��p�[F�m�{���rpxb�F�J�v��Ү
���S{� ��O�s3ѭ�R]=��z�櫁��TzƂxZ?);��^���Ն\	C-wq�2ф�>��J��-�g�` ���E�)E�iF�)`�GĔ��9�ln�@=�R��6軪-la����y�i�tF�&���|ș����ӣMm\ܙP��%A�b�����o��<���o"���_�z�����M���$�O)�Dr}ev{�y��#�p�<���Lv���7)��B|��kk��a�����Cs(SF�HpI+�N�
,�'���sk��-�b/#U��p� OEdw8x���AD���^(R`i�}�����$�5�$l�o��E���yC�Z��h �زM��P;��t*J�3Bs�
m*5�9�6`��-�0��y���Q��M0J[;Dh�K3���A��BJ���A ��[�7��/��-��3�JHm�R!d��J�P��p IĠ����Dy��Ӄ<�Uп���+�a����8�B�>m�~��%t�!-.�jQl3� "�hW�`��|d��U�YS�r�6�^F2|�ؤY,�yy�x?�b6��ɇ��f �Q7r	Dt��@��m��Q2��5�4VE������m�� �y/��)�J.o��ۈv$���h1�3��FW�[s������a}k83��jU���츦�8����� �GR��z0S������i�q�5!������_�&2���\I^)T�uO/CM.��_�R||p��$	5�MfL>8,`Rq.C�l�%�V=��+�-W>��
�?�kא�$�5�}Sp�ȫ�&"��dص�ux�Oj$����tmі�`ߧK�{�>���CT4���Ы u��UdK�ȯ(�����҃V}��r$=�N�A�!=T^�+��%�dt����x>_�6+�(�)G}���2,���|�E|���d��\ְ���S{)^���H4o����t�U�KȚߺ��X[��-�+�Ivl:B2�H���=�L�R�i��&�w�N�'1㵝�9~G�l2 �t6�d{��rg�#��D[��S��k�}��u�7�^h���i�P���#�}��W%���Wи��U�v�ܱA�&<�%����c��VGy>�2�vH"�[��!$U_���Ӕ��A�7�2�0e��0���Z␻���(�>�d�9RH��ky˨�+@�/j�/mw 5�2��P��v�Lʔ)Qٵ� z�.�3 4E�b8ZG��h�aa�=W�H�T���
��ެN$qeh�\��ݻ|�����cɸ
�Q��*�JB-�n�L�j;����F90#���{�~�<���XՕ6X��w���N�5A��닥A��љP������ᆤ�i6O�e�ǿ^��t�i�+�7���L�c���S��9UD�b2�,qi.���C/>gq���لJ<�R�Z��#�ۦ����ɶ������aus�;����v��_��LYd� �̻���̼_j�EJ&6���&�!�!v��i��a��˹���+Qr&�d9t'f�Z��g�PUf��6b�bYm� �0o�?A�������fǋC�}06�������Iu�ZAGk�])�n�s}3�T�"9�ҏC�s�{H�Ȕ%�6���ö�3&���a	YI7�^#�mNQ��o@���la$��.o{~��}�Gv>Sy��
;���	7wj�X`����TdǛ���`dz�/���7�)�h�B%AFUo"�!8���[0��Kc�d0�X8��i3 �w����S��뚟��/���g4a=�� ~q:�
T�!���9C���T@J��"h��h/�p���YQ� '�;��@.���hw��JA�*��jm�����&�28���k:�G�>�����* H�j����Ɖ;���TQ��^|��|�n�\�f:�EaH���#R�#��� �V�H;y�~���p:&�W|�J�FhÉ��o;uɒ�L0 믑K��B&:��V�.ڽ\�����m���1�֥ �t�U��)��,��D$��Xt{��W���U����>ΊP�|�}�Qw�n�&�N�o���;�P�u��McTh�b.�����L�����xM�/g�'E(�Gs��ae�uHb�S������̃&T}E4ً�����U�bM�5��"$���-�;�&���>�������YW���m@���OFx,z6 :���%,l�����&[�c�ƾ#�l=��~����F����!��f����	'jW~�����5��+tG$l�HoXd�v�~����Y�`���1p9jv�	s1UM��H����.��H�u�HW6/vq��P$�Q��j����7/�-��w���ikF�#7��68��^�xW�6l��C�J-�wˀ�-��c?o�WRR��R��Zf2�C��=�.7>����w�!���,
�w�O�V��(�ꏗY�\9[�<��aaFHԜ�կs]sW�o{0?����(����Q� ��ϰf�M�ㅩ��<��6���%�ݽ��X�<�6��L�G�v����y:gg�����C��tPT��cB�H����F��WݿH����GyS��<��zڋ_���zY�lԇ��"Vބ-�nOH�<�t�X%���u��ִ��0�F,��"��R}�^{�s�&Ѹ�,�l)|�n|iH>���JhH���0�v�QU����%��L�����#��qT�R���G�)S���%0�a��~zmaaW��;�L�Wc ���(y���'C��ST����WE֬��ց5�v��pq����b>T	!�ۤ�s?G�CNka-������a�S�M���!iԌ:գ�J!S=�9=�f.��xR�w��:�+A���}�;�o�R��o��=9��l���f��O��](=��BŒ�L�0H�FE"��̑s�'N]��/�P�\D�PV�����VD����d��m�(X���D������yqVQrIX޺!��R�$U�ˈ�mG����h�h�Q�=�ۭ�wLx� �$Q�-��M�����qQ�3���-�i���Ni�B OC5 	�6%��m�|��f&ڮ�8b�b3�Xs�*�4s����pր�
yu����w�C�?��[9��B����M�f����Ja�+��j�b�:c'w�Lm~�I$�l�'��tn���c�q�7aVᢺ�fx��O��iP�Vm��j��v�k�����6��� ��q�A��gT' �����io��ڼ�aN�Rq�A��T�g6'G�����x�����E�����
���o��ÓMV�KZy`S%dzf�A�y~�	���>���+��{�ȠI�ɚn����YJ�k�?)/��a�dr�<� �u�^*
�T��V�7�Ajo�����"�k���!�=�4o;����߉���c��*���QC}�O��Ň`�A]�Ц�)���7��u� ���F��[wt�X
���96x��+��]lś��u�Ľn<���,�(7�
�ٶ�<�$�bL@��
IE ���ˢ�>�M�G 28��4B���P|R��L��C�g�*hȅ�Fӷ��J�ɴ���z��|aOm�7�Ж/���uR��}8�"*�|������Dx���o��BD�Cw���0d9Jb������{��Y3�y��6J������|+S>vo��'���^7~.e�d�}���\¢��2@��⓫���}�]�6(�|�{W�ݙ0��ͣ��;��^%���aˏi�v���\�v뾴*<Ш���̝lXY�YaK-�X��!nRUFg@v ���LAah�ˢ�-�+{���P(e�c�<�F�taY��8m������ �\I{���9߲r�W ����B��o/�hg�~-�ɿ6a:�A܄B&JhM~�� ��Y]Zۥ�ۏ����j%z^�ߗ������P�]�� T��%��g��h�}Խ�9���hH��˥c��VlIf�Q��ɘv8`W�1���&�e�&R��^��6���U�8U�p�wY"��]#���4�@� ����lHy�ն4󇞁`H�e^��ҍTzR��FF���Is�w��� s&�	!��0�,O�R�XquA���L"3�ئ/��5��G>�������P������#B��؅R�4x����k�:�R�������Y�DEn�j�&DcSs�1�B�:i��������б��F���l�N9-)Z ����K����ؖ5%�D"D��^:CzK])7\Ⱦ�1�Y}����dE�`�w[�p	�������5W�b�^�i����΃\in7��|V�T	A��(�-����hɒ1[�r5� 5�4d����s�8s����6C��|�<�����v;I�#J�1#B$�_�T9)D�Ӂr��b�@�C�?C�p2Y���������JMEu�mA ,�.��]U2"b;����_�����d���JWʣ�O5
c5���:����}�3[9�2�@�-���(������-��:���-o�)��8��x~���r�7)k˟!�bn:��&_���S�z��d�E���;6Î��b�{��{�<7$�?�M5��~᤿�:�S��$�!p�a�L�=��SJ�Mt�[s�[6IK
����mW�GԘ��	S�`�`�7��6��Q�����7 F�ǽ2[~sTb�P�Ui5�`{$��2�����jT�߆(����^s~O�� �'=9#7H?r���s�x�B��t#*�'��"����qc(��w67"�c��
���n�a�Xl.ĹJ�]��y	E��4kG��R��~�P8I?��e�O��(��&z/�U0�T�=�HVr6z5�Yҳ�,��7j��XX�	Ed�� �L�j����1�V7����σ�ZDV�^�nOn�-n�03}g�� �� j��gl�T�T��,�w����e�5�~Bj�����$��p��[r�=���;���V�d�?�p	Ǩ����_��XQE&H�	��4ƌ�v�x"2�;G�l�a��X�e�xH��9����7-6Bv�b��χ�	m�se�|���0��Cvn�냪��2��*��/�"1q���Z�xg����ذ|�FE�rt����F�BJ���O��1H1�>����g����dVgw�A����Wg��\$]�&��NDE�+E<T}5D؉�G�N��i�7�YS��q ���O�G��s�f���L��]+>r'��~Ԋ����ʲ���&^��)P�-���%��}�����?G8�i�hUW6%��p�B
�cHa����*ʎ�"6�MU�U��Ij�y��6BcgP7��>�䈌�0w��m���~�ا(�j�ԅg��!�\;�<::�ȽwaF�/�$�����_W�Fm��{�j��d�W�<t�E��ȝY�z�l��sf�iڴZ|�N�W����<���i��w��)�K���)��0+���[bm���Z�BE6����_|�O(a۪S��ն&�B2"M��;��:�Uc�R��\�A�hE= BV��_jX��h��9$ �ūTq{�x��ȩ1*��-N(���,')V���]&�W�p�\�굗H�M6B�m�(�=l���s�ZI�;�x}
�,*2uʵS�/��D��_"��#�����Un�1|�g�V$k���\
A������yvV�����u$��RJ>A ͇^�o�m|Ԁ�bU�hrY)�p��J�M�tHZVM1���P�0�nm
ըA������чroUj���8���=��t�䵧�@lZ��9���"�<\�S&&oG�<���4�s�U[b'H�K~4ެtEl�ˎWE3�%J���8�{)$ٶs�`Xt�l/+�Bҥ9G�����#��߰ث��k��oL���Vo��pjʚ��V&TIwH5�����R\Q3�J��}E��V��38٪؉=Ѹ�Uh[�z�$o�w��o��`w��.Z	�Һ\��Z�y�^�dq��x�2C���+�)�8\+�[�N�Ǩd c򎰨d�4	����#�^1�μ�\�e/�q�4P��_;n XlP�%ҩ�g ����'�&�5��1�n�t�����S=�U�ǳLQ>����ԡ��Qa�q =k���OVYt�班8"�F��茡��Ivyx���/��bϭӆ�p���0��=��p}�(b&'���b@up��j¾��\�.�Ň�3I����c�r�8#i?R��w�w��W��8�?5=L�<����lP�y.,,��%�|�8�9��W�{k!j�ێ�EJ��SI�96����"ۃ��A�{qb���=��%سT�f�m�u䈎��Z��_�K�|įC+�m��W�󼽏�K�n��$(S[珤��c,�IpP��mX�����4��������G�N�$�Fnk����B�M��O��@ƕ���X8KAw���z������D!
t��Q��֮�
BRBLL��y�b��A�<v4E/���	""��1	7g�%zxH�u�t�^g�+k^���޻o�N�9S-n,�_|�mm�&����^�DB�T&'�wX�����9J��h�	���{��8V��)��$�⩘��N�_�K���*�I]Z��ӎKR��=�:��U���e���i<o����� �%�C@���qJd2_�pĴ'/i6:u�ɧ������Ĩ�ư��B��H��l��f�U Үͦg�.���B?bƆ�=�{�""����b�-��Z��_����16k�j�9�c��D\W��1���vW��咽�-�kN3�!���2|�;uN�Mi��K�Z�]���I��}�_:����2;�Ǩb[��i�9��� �T�����)֌�o�E��Y��2Sr�Qd^�����T޲8�����1��%�ݒ����T?,�#Q�p�#;�ZAF�O���#T��</ʌ˙�ɛ�%��/�1��l������z��=�Է� �OM̪���J����o�˷�..=q��b�hq����?�^.�N?��"���?��'n<c����I�]R���x]y����Gܰ��2����Ner��D�8��F�F�v�\Fi澳���Ջ~�:"A��2�&h�cA�"���B����uܙJi�"���2N�x6n3�$\5[�V�>r�ё=�p���w�n�+Ǫ�||���4�v��5�i�3��م_�������4c�������}���e����<񺠖4��G����%�>�
��h��3��?h�/e�y��W�'ʛ����sm�%M�1Bu�/�XQ�q] wnW�w��[
�IČ@=y�"�a�7.��I�l��~骰E9FC�&��*�I�lu�j���{<����v��äI�!f?%����q�_�*a&���"���S��2�T���t�s�����аj��CӠ9��<\���0|��>,�Qf� ݠ�s3ﳟ�R-�;{)M?b��c�(�/�3��ٽ��d�/hte؂���|txw[��f%�� C��Ta^�R�Aj �Jm�M̬�o2�	��M�0��-��=9��]�����ҁ�^���O$jH�ǘىK٤�j��"]$�/���n�%MY��'�=L'�䓏�s��K��Q�{X���`b�dY�y�9)�~CGᛷc!B�
8��X�]�Avv�$�~Q�X
���E�.A��A�������%��4z�`i7P!��@��J�E�����S��3W����I���&�%�z4�L�Ī�\u��S�~��C T�4#��%}��p��Z)�[�Ճ�Ex��4L%f�i����I�f���'`�w���SK��|Zis�k�~��7� 	�7�Xpb����Ce�X{�b8m,T�|�n5j��x�ݪ!�0��� ZZ����~?���T����U�x���v �������=���;�ãޅ�z"S�o� �xĮN��s#>�]y�\$߱����$�x�^�3��e�8�D���I��GI&�;~�Z���N�МϏ��	1?�"�<d���*l,x�T��0(�9�3��B�t������A�	\����T-_q2���r-�.�������B�n[)�T(��/�o�'��9�%���߇=�ٱ���9�l:ެT��Ƚt�0JR�_\j�R�E��v��FSݎS��E�v�~L�'�LJ�Y�8!M�s�*K(�ph��/�p�Pvw�1O����YdE��i$m^�Eb<���
�Y�����Q�n߮D���ڶ�Y@8|����5�he鸁.�f�y%^VC;E�6d�?��4#Ni�m��,]���E٩7R��=�UZ3��p���ΠD�����	�'�})�v�~��YDY@��׬\�����op55�x�Pܰ�M����[󱁢��X��kLCѣ]ĭ��8�C/ɕ�_�T�dj��i��+�� ?��l0}od��L6���5�%f�U�[=�&q=�h/�����Ҙ�)l4��t��3+�u��(z#"���@ t��5Me�JgB%v����H�39�]��A����k��~����ΙлИG�u��4����B¢	{���M�(�IA+�mo�`cm;p rfZ",{կ�L^����%�-���W$�����kl0hg`��?�3����>�4C:B�"��տ�=��i��g�V����E�v�b&����j1āLpIq�m!�*$*���#��~m��3���D�=O��;�\>G�3�5�$aD�T���<�^J�U�q'JևZ
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@��[�nL�v�Q���<���Dxv[Gt��I����c_ypO��gE��*R&5��y�0�8l�6�hβ�r(�aI >��>������P���S�(�=]%��튇R�����/��-��^f�d��"��묲38\$j�֬h�f��d~H��������c�*A{�|P�d�W�A�3���v7��L����Z����lb�bq�����%�y�y�5߀�T�ixl�Ѝ~9�|Ͽ��~�|�IoN�l��_l��"V������O�Jd��pIMv3�:A��~� 7:�Z��7.�m����,p�D,j�Y�.�d�@*~Zy��!��ݡA���������fW�3$�.��`��/��\S��:L1�d���ag�:��
[A�)X�!+�-��g2�y�YjQez�v�.Ӳ�I�2}��D9Ky*>_�W_m��-��?��"���%'^���\��>�8��gk}
U�B�vK�_���"�O���$?�7�D0-�Zw�jf<%���w6Z��zE�������϶�6�x�ܐ{y�,�._� 6��|��l�� TH&��{ۡ��	j�ཥ]�P�w�A��/w�����`ј~�Q����_��n:�9����otZZYz@���SL�"�⣌�[�0\'[��6���2�N��^dX�J��z�[��.��x���RI}Ɨ�U��-Յ�ȱ�	n������Ÿ�3u�@N�KtQr�V7ѕ�|��c�x�?�qD�+�Ŕ�����������Ќ�o�ʳ�ߛ�@��n�.���}�^�#�(FQ6烔tld��{��y~�� �u�'u����ǿ�O������������^�rf@�kg��z?dE��
ӵ��{Y�®2t_�[�K�U1�.�"�lUh��;Ю^<9�Z����T�^|uhw㪵Lѣu|����������P�[~{_?pf}�	��$����CVB?��n�^���������3Hq�c�:Ż���^!��-㼍r�9w)<H�Rb�/5hX�a���wV�M����|������E����8�xv��<Z$�t�Yt @�H�����Nȟ�P�rc,p>r ��{�X�"o�S�q�I2#���}+d��|n:I�Wh��������GR�D�޾�썺�Ǻ�������# =�あ���Y���D���$\ 4�`�N�@u�V�a.tns�1�����}߼�}mϳL�c�X��$L���1���L��k5��T��@Ь
j����/N���mb��P�����ִ3�ӹ�C�4�b��0���,k��[	hQ29n�\�%�s�>�ᦦ��̊��8%軼Pvn�"t�����B�<���<�BA��� ��ح�bU�ڸ��b;�jK��o�m@[7"�h�n1�	l�룶XwY�:��{7��:���}�"�>r��2$C^p� ���2��i��9��I�ge�H��Y �}ю�G^���� @l8�5�i�����mu,RO��h-�x���W��s�yףߓt�y A���/+u����Ha�z��է�ҕ+�b�S!�V|�O샨_(�V�w����º}��n2z��D,|X�~|����o_м�H1T��P�� ��ώb`��ø��9��ː6!c�r ' B�[F+��(�#�"`I���4	�M��@4RM����l�-����5,�TD]iQSl�ޚ+�����
������!p�Q��BV��I����%���h|�v����}�p��^�:뵦́�hU����/�ՠ%u��~ה��t�ץ	Z�%(p����S�°�@O&�m��b�&�mΆ�ֳ
�
C��A��cc_���A�����K��w=��_�� .qCzu���@Ҩ��ɕo�B���V[��O�(�2+u�t��
�lݶw6�G'�-ѲO_Ƿ2S�i.)�I@a(&�׌j�~n�������Ҽ��P�7Sͻj�L��>���~}*�n�@Gf�X�!i�������������R6�$�{ �bI�/q�a2�$���U�˯:h��t�C�E�ʠB�7�!��L�I ђ���Y�gpi��'�Bѩ~6
X�}Iy�kg�*�����5ԗ4!�:����,:8�j�:A�0��J\�q��$�@�	��!�+��B��J!{*%�)��i��^jx$��hM�(""i�KS�_�P��V?ҽ��3�K�����>L��
s4�S�~�[�7k��]ec��F�qRڪs��$6�lх�DG�W
S�v��>�vpA)1�^=M1���2�`�k�{TB���^��ӌ4��� �{�E�,1���yb5H�z-
�&p?�iK#vC���o&��
{��k�D����v�87$?��V��r>>Il{��oB!�h<�`�=��3�C�)�f	�/L4W�!H�Ex���=����kdT����O��k0�C�	���W�R.4H�Q7��mp��Ϧ�� �KW��@�t����LBb{��C����]��2��#�R1�-��ź�;i?�+�"�Ō�Ȥ��9~��ȫG
���
������ޒD6���+�;3������t��M�+6���`�����^�E���n��,��SЪ84AsZC1�C�ܻ3 ���0T��f�E���e����r���4Ή+胏��WTa���j��h-f��[�	]�X��n\�L�E�@��(�:Jq0���&��4Z�*s�X�4���G�'�P�S!E�������W�S�V����<'��7�{ ����ήdg8���)?��
|�^���*����3ш��4�;�Wķ��dEԮ�^i���0�q���B�%�!����$��N�9�G���������G�w0�7M��U��_
��,gA0� �g,���rh�b��F�S��"?N��:�gT�x-�M�+4J4�uw	��^�J����ۖ$�fpw�����_ʵݮ��\���+�$-f[!�ǎ¦9���� �@i�&��Q�=�\?�\$�i�
���:<����d~����+e�D���NK1�,i� ?(�-%D-��׾����a*u��]��Ӆ_��I%�w���g��=x�9���vAe7��s��% @x��w��z�Nq��s�pb��U���3u%H�z��:'۳�m%��C�%�?�������?�K̎���>�U�v���W�A�v�wSrU%�
K���l"n�K�gq�T��XC�{���u
�R|*]7��v.�ĝ��f������R:�[�M�)(W�9���3ee��	>2���;�k4''�t$�Yt@%u�� ��
��`'+���h�*|3k��>���0�+U������I��Zgk6G]�r�U�T���d��u6r���}���84�/�V(�O2�IU�K*묕��nN{"�g�0_����pBo=+1D�3@Ԗfu/P�;�yf������uW��g��p�e�]�JA�_�v�	 &�=��9* 7t)��`����^�~;"
�I�~D�Đ�^�FE����EZ��� 7����
�:ȏ�V��j��C�mx�U,�Z����j�)D���LF!�m��5� ��Y�f��.��C���[HA�(���y��3Q�Fb�re�����?L��Bt���?�z��$W�u�0ʼ��Y���SeG=U�:�n�(R�]��l�ڔb�0t���nӲ{�h6>��'���U���XԱ�
�n�]t��4:��n�LuTN?L[(`1*�����	Gw�p�]+kI�'氞'�����Yi�k��@@=��z$���g/�Lƛ���̄���q61�-��2��� {�+̝x�$��B �вHxM"U���	��>��[,o�Ѳ���$yY���6?�^ޠ�n'd�.[�>�^	���FXg���Wnc�:� <E\Fp}TD��}�_�s+�y;��t�������uT� 3qV\�<���&�$*�=]�9�GN��:�ȫjAW�n�,��^E�1�Y7�5v;��T����Ξ��"9r"R���.�|�0gˀ�8��D�$�����a<�ja�����:�o���{Ǆ�ʙ��f�ٍ�q��%�@��{�0��U^�j�޷|��������ٴ�|�}���	�����k�0�"�K����@��o������
�*A��FY �f	
g@ѷ[�������=m��V�g�W�tIɂj�����B
̇���"�_�D�����B��j�	�YQ��X��X4����RK�;)Bc���T�u�ο��r��F��KL|`�n�2�/��\hL��-�Ǚ=��1^Ƅ窿��M+�<i28M|v�ŗ�����ٲ�z?)�C���bZEx��C,^�-��eR��Rڌ�V�e?R&��"�:wj�d�h��@V^0�?�������}��w�-c���s���?^q�fi���L����Tm�)�91(` �2I���ݠ����:���P/�aU�F	J�:�e����;Q>���Q�͂�k� ����� L<��W .��cM��04��f�)4b�W%xk!��c�gHA���&�� ���o x$�V�ʵߌ�F�O�mI��㸿&Xh��૘`f/���G�xn��d��\9�蔫4�n9��.�,�D��Ϛ[�i�*/�fP��+�~F�w�hl�"�^T��ު�ꗿ��.�0	c74D��ip�lB�U���ߜ���i����?�,+vL�$p�	��l����C9�H���\�ښyg�Y@e&9�|�Z<Q��(�E��:
���t�,o&T��T����fy�3uA<d��!��dwڴ����d2�fC���9���Nq�lp��Z��$B,7�쎔��R~�⩘�_"M(�9$5��>�^�voO��d�4�#k3��l�-Yd�V��dC�wFK�W5�9��9f�G-��'N����_� t�;�'����F���~���R�f1ѿ�������'�hm��Δ�l��#�@	�B6���?
\�0�~���׿�
���*���D)o>dsb�/�>���Ǔ���K�:s�M���'MGo�Z�>��ds���b�N�u=���ωy����Gs>��?����ޠ��H=���S�X2n��!F| �	f�j��5O8	%�/y:4�/Y�$��탢��ns�R(�
C/UrƇ����a�la�r�К���W)�7�/�B�����8�准��?�$W���SuU}���s�ְ���b#h�0��p�������a��h5S� .�p���\��B ��KhX2���4"?���8 E� �����4�q�>�%I��a�y��:�u)�w���<�e�X�7_J8t�&��b<`k�`��T�|S?ǘڳ��Ȼa���~h�"@"R����R����.vqYِt�Y�tn��5�[�|����*��H�s��R����s,�DV�ܴ��y�5�~�_��!(�2�,!���~��w�	��-v9J]�(�۴!X�v��D�/���*/��
�+� �Kƚ�ɲ0��̫��]'O�V+ѨĿ(��x���	쇵#� t�ۗ�=$����.��"�~�;�~�%�f́���4�M&la���s��2����8���E�d���[��N��__�/���W	5�!(��U�3z晓cq.�g"SS���h	� f����8Nm�9:L��#�ݬ�"3WΫV��Ʉ��)��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J ��PNm�z��Q�o�� �A�k�@����ehh0�_�Й�ŏ���r���' �7	�1��E�j�l�p<��)�Q�t ����調;�,�	U;|���=����v^Cg�pI8�~��1��C�{HI��5|��2!��B�$��h�:o��
��]V��$9��#����'�R�U��_�A�@7&Z����N+�C�d]6��σ�y$S�b�8;0<�60���F�x�yO��/I%�h�a�0��� �h-@�Ч �v.�o���ٜ�����ʌ�'PV�1[�bj�|\~�����E�r��M�}���8P����"�a7��Ƨ0<���ީ(8��j��x6�����>�G�!zZD�o�6�ˤ)��uV��\C�S/"@���K����o�?��m��+�X[��Չ�9�|��}u/��%���냡ш����DIF;�D��`�S�Q'E݉�EJ*��οt[_zp��X(GO�����1H��Qa_Y4�K-�C���X�Ѹf��;����9v������n��Q����_��3E/�Π����œo
̝��`�I0�o�V�j�R4�gj-oF<͟�&Eu�$�_���X/��Y�Z���~�;��3��h���F�.��H�7�0(����ȫz���J��Dr�Ӹ��� �`lms1��Z����z*V ���1]�*%�&SEDH[k\��'����5z��]M���g�r�w��Q��? �)��j�N�7�Z[L0<�w����d��h2�v����&}i'�*�%7��2�z�)7!D�������Rd��:����E)!��?L�0Ĭ�Js�y����uC�<f��:�+UlA,H��$��������D5��g��PY䃿dB�F��ɬ�o͔q�sQb]F�I�>Z�4� �h�|��s���Q��4a�l �ְVZ�ȴ�],���
;��WY�\8�J�������GpZ��&�y1���]=�B�� �aB�V����~�S�ů���EK�����/�bd�6�q$Bd5��c�˫�w���,Z}OMX�4U5��4c�ڔ=4�������m��l�NV�f7;�(��#�*-��"�
�T�q�h�(-���ҏ��V��-���@����A� Q��I�� H7yt�u�p��L��	��E��œ�ĘC>��BE�U���*�"���V��.�#���滞6�An�Y7C���1d��yh|�͌� �QpcX?y���#�Y�5���|L��ɕ�-�ĭ�����y{N��z��F�x����n����6�����[߫c�:Q��4(0��R��fu���vMB�����$x�Y�sPn��_�J���ZJ�sx�����9Uj(�
^i�7���x��gyx�Z��������]�Tw���䮕�� ��ܜ��% 
S������^���qc��4��d�c&Q��ֽ �?e����Ѻ��Zz����N	l�{�����������
�8֖:��ߘ%�Z�����s�cZO��
�p��_N��GA+y�ٽz������9G����@��a�+UF���h����/3�����~�1Í�<��Q,Q�+�TĊ���d�����߯]rx�_t%�Y�������P�����w& ꃻQ
j�VGE��kT>z�[E2�]j)��o�� �6�:sк����6���:;Z�����VPkN�/��S���/�-�7HI'En{����� N��!����_��A�W��%r#�!�IG0Hs���m�{�\�-�c)�r9�s�:m�H*/e��1�Z ��8KƓ?�	���lV}`H����tZڠ7���/��Wj�Tj �{O�Oe��"<M�'�W�A>�+�I��"zU�g�6�Gp`���?uݘ��ҷH������vO	A�Z^+�#{;�����[=�Œ���+�Y������~h��~�nֳ��v��Q�u����,�ێ~��8��1BQA������L��-�e=���&n殐1�?�,G�ۛd�����Cf�c����+�]�}w��¾"SI[��3ܖy��6s�rY!  �o����uB�N�R��G��wE���B�������ڷ��;6]#�Ǉ�E��1+��XF�q�̇��~k�`z�`�ۻ��h40�Uz��쉿��J�RV6j>.(S�7x��" �j�И&�S1��Ԍ����b�	��Ч��ל��b�Z�[��;�N�!J�g�'�@�\X��Z�P����'��ti\���+uo�y��*�������O �{�����OSEiz>cHq�
�t�׭Sk~��e�h�\X�;:��v�/�_�¹�h1 ��S,c<�#�.m�&�PmZg��K�@�za"'�$�P�.ge�o�He���[u��~�UM�r� �Q^�����+ekH� ��!aŽ>6`D���w���6`��X�ͤ�r�ǝͅ�4 `�<�tS���{�ܵ�$�y1�q�`Ɓ���D��Ez���]�{�`���;���}t8������LbY4�c���}�����?��ͮ����	�� �@�)߫d������ʴ,����V��2�f��A��*8���S8t�磊n&Ӷ�'�T�,�@r9�uS%�@�=�qd���� j��s�Y	(޽�a��
�N��G��}��I��GP��cm������Gt���̥��doV���\���TS��+m[O�K���Z��'#Q��_��w���	�b�f�T��*�9���98��5Q��Y��#��F#tϢ+�y&���p�#�sU	�1�T�I�;'�I�.�H�8Ϸ[��I��:3TK�\@l!�X�B��!�&��w�W�,	ҳ�h�uK(q��r�l�IW�:J8�L��?��W�U�"�T�J���
ǻ��;�Vs�IAd=%�Ez�������!�\�Y�rqG�K-��l Bx.k����2�R|xz�;��9�� ��w���2�������pn|��¿��gN2U��~�3�PEw~k�jv�^׼��JY�VX���!�tlě�L2�p�l	N���Aik�f �mg���X ��-�BO{�?7���:��ۙ$��	)�z�S��$3��Z4hef��&���:q+�"��cj�����v�ObŞ���.��c��w��G3t�N���?*E�G�2tՁ:���z���PO����%i�K��w�����SЈ`r�u�!\���@�W��֎,�60u�}�js2PK��m*y$���W�v���BL���;��>���N� �"Ht�|)�C�6"W81r��C�{��gST�8�\��.x�($�4m�i��]�xTz63�h��$p��iby�-�pE�oc�?R��-
j��No8R�ny[c��*X�����X ��O!�G�r��Ǆ)�����V��U���&
G�N�BZ�"c^�f��7�s�L	r��t�)�vV�Hm写[��I&�	�eF:��T	I�00:^A>�/}�ѣ�`�k�K7d��ْ�HE���`�b�z��g!㵝A�����ٱ���>A#K@Ǹ�s{g,�$���E��W\\c������ mR�I��u�x�9�T�t��Q�{�>v�[m���"G�&Ƀ9�qsh��L��fU:N�Y��g@��w�nR\���̈́�Ni!�r|�a")\���2����※�}2���/�cۤlt�f�Yz4���'Z�Ç����cm�;X�<?Uuu�@�2�ؙ�v��й�y�k�^����Y�T����@ư���^�M�ny��Ky�b��;�8���x!%(^b*�����Z*�`��(T1r�4^�:d�V`~�'3s�i�68�x��pj�A��a>F�u�ԡ�Edp�k&o���"A��NV��s�ƭPj����ʚ�ʏ��F�� ޽Q��C�Zh�2
0�J۵������\�����^�[�i���Wڵ!} �` Iy����$ Ȋ���1��'4�dIӯ���j�ܚըzCof�oF��݃�E��R0��w�� V} ���wH"�6�Nx��w�V(eF�zh~��A�}9G�ˀ�4;��������n�k��3�"�ֿA�+��&����̫����л���l���M��gX�=3�=|
˛I�Փr���������ݐ:�2�����)��<�XN��.R�����%K-��N�j��H_p��Q�Ar/g�
{z�8�)t	]�����M�9ҽ��������/�Ͻ��aq�&Ts~S��x�M~�<H*�|c6w�����Џ_L�k�"_\�r����¥&�������j�Ф]��'�K׃�;��a�� \P�Z�#+�g-����f�E�8�Cš�gq�1xEԒ�`�Hɐ����֣{;�����Z�)8�����eC�Vc���U��R��Qwֳ,
/\ �����Ơ�h2��Y��~�<�~&�I�b�W�F���N7�Ǔ�R��p<U�0����a�\gw*^�n��T���*X����Զ��:��>U�O#ʤ���`9���u�Y"
��R��S�c*���	�9-TK��$o� ���M�^ȾL���e�^�f�ˬ{��DV.��d��5�O)�%�BRb�Ce%#;G;�t~�_��:��T��)t�mP����K}�F�m^�_'��4\�0�#1�ޛM�D��
fv����y�c�:�|6��7ʫ�+mG��J,)5�V��@�l]�2 ��$�"��$�oLo;P���"��.��qlS{T�ٜv,�'����[��U,���S#�G~y��Ԕg�,m�)N���Y�je�������ő�M~������,"��ޤi4���;�g���!���lPݝ�
'�g*��=��?|v�d�
��M=!e
W����@�K9�^+����$G�Y�7�&�E��y�:�Q�?��_�gM�ƶ\i��rS/����(�zv7f�׾v�Z�z�Y�rn�I�o͑���ޜR"����� $�'���6Q8�$��s�r�����Ȥ�G��A_$��2o��l���,EE�/�ܤ�ӑU�t��]N�*D���( 3f�-�Rԫ~k��"3tء�º�~��Cө鷧��<��YIT�y�GZ�'���|�Y�z�/jiZA�Yq��o����fXX�d��F�8�T��W�*l%/�d���*)L4�jY�&{��(���c�]<���}:�p���ܧy�{�xH�vϪۊŶR�Z�zk���6�jgqɐgc^���ZI���&&����/����P1�{H�lQgh�����H�u>:uC�A�Ҍ3�oؒF����ϘV��㕖FƔ��j%VÙ���\���Y���n����3/2㍢/[<=,��Ja(�AIh<=���(E��<���^]�p��=] f���ߝ\�A�r�Ӓda�=S�/����g|=������|��7����������e��|o ;[�,�ݬ�W���+;�6Ԃ�xZ�a�����&���pI�TϦ��[����OE�����b/e���[�Ҳ�`���?p \�M?^��pC��%�� ~~� �	ei�_.y�7j��w	V�KZ���4�!S�f��d�3nL�yr���n����4�r��,�qBU��]�+�=ka�<i@4)nQ��XQg(�K���sm�ZT4�=�y82�MoT$��f'hG̜��M�6Y?����n����uڛ`�k<��7C�v_���d0<\��p��Mj$%
/in�p��֨?6�⅊T9�G�,ȥs�ܟҨ��-��xM)������|s�Ma��C�i݊F�*�����^��a�l:���4fma����K�Pl�{v�����R�Y�r���nR`�K���#�.���� ����Jpn�4&.4�-�S*�J-�*|]����d���¯�h�b��FLO\-r\A�k���@<8}0�
�[Y�[I� �4x ��X�͖#�*�yj_������RHȖ�����5�Q+�t��Hv|���Ɋ�aK>�Z[~�*Q=�`SԬ���k��J����J�����S��'*��0v�-5�BA��#�Z0W�$+��ka��q˯	Br��H���r}�U2e�������� v�c�b��1u���o	�L&"���Ħg���s&��&b���叾�ˣ��@_��΀�j�nϪ+G
�4�ry#o����Qѽ������c�J���m�?̙��>�����cM�eU��'������5�T�
�\������^���}�Hx*+�Ƕe��o]�_���<�I��{8P�����4���'�с�m}�i�@>�,s_�g�!E��1/�gl�1	T@����`o�z#f�ɮ�*4���w5�������j#B%�ЖA��8�Go9M��fu��! ��3�b�ab�����!ْ
�{;�Ht�1�.:/:��V5Ed9�er��r��5�h��nh� c�C۩.�uZsa�(�5/a�KVI�iJ�=�Xܚ���8�7r9����ޒ�g�<o� 0����0�"����w�4	3{p�pԆ�xd�<��{B��ړ��`ڊ}��,�j���-f{�����@��b�n�y
��O�wib��2�D�F:��)Z����:Y�j�S�jW�S�����װ��:�0���=���ϭY�lRkД�h����{L$%ܒ_�s�]|�3��ɻ*Ӫ�90{(M��T���Ӄ*�9�]�4ʑ�S��&K��`���.k�d�#�
�d��(�gW��y0�Z[�$���
&�c0�%;�V8�zDsv+�ֻN-�F�܉U@��ZUBn��?��ДЫr��]��L0~�)�-�q�X��sӰX�wn,֖w�A���*��V2������	�`tA����rg0��d,��O��Xx`���b�s���O8������x�x���_J��2Ϩ��-\'�Yi{�
�}�fd�����5�R
�QM�D�2��֤t�rt��K?�^h�%S'���K�h�!�윸T?u���d�I��&�1��5�W\t��\��Ƿ�s�H���%�d�3�5�L���_�����_��ˋb�5ߵ�9s���� ��(6�%X4g��5	D���s�Q���+��k���E�P�pH�;ȃ~_�$1�.�C�<OÎ�\��m�i塐�����l��h�ZVȇN��g����͉pU��x`��r�8ſ���H/m�v�<����0ĲWn�����-7�ڣ~�Z+�� ���}*H	G�y#ݞ��$�Y�R�'ݼܻ�2[�?�(����An�ЉHb�]j�*��X���S!vh*g�Zoܚ+SVCdT�(X�5X�AఫȱS�$��Z(?�������K[zU�U��$�*+�3n1��-� 1L���8b�N��w'R�|g<K~ܔ�親~4����9:\Y�7�ho��Z�S�c�Y�SS��$j�8�*�dp+/c����F���"Y�黍Mb�D-�c���y_) �۳�����X;J�r���� �o����>�-�T
^5�0|a�Ƽ�]�׊�o�KT�x��iz"eE|��w�����
fg��Ye�A��#aLYk�1��/y�չ���?�_q΍C|�V��/��ݙ��i�FC=g}��aM�K�,7����ɤ���X@������8�����QLO�Ge$��ɽ��?l f�����#�y'���C��vQl���//l�A�prQ&��"ފ*�k[�g����M��$v��W���}K�u�ʯP5n����=嵿8!+�*���Q}��xue��2]����D�
���|�@P���PC��3�F��䡃����',�k�3��:./|�PY1b�����j��$>Sa��|�f:�x+ ~Ԡ�7���E���>��׎LVZ�^h�:����/�L��X ��,*}�(���/�G��8���W��+M_sT���|�fpʹ�����C�����z�W�Yh��I�N]��S]���SW� �Q#`����M߄[q>��.$�J��/I2�<����]2�Ɨn�WA�ˊpM�PTHReu�����k�]�Zr<A��{,D�O����/�w-\ X�yz2�M��87�3�)-g�D�7��5�&�c���Y&�F��J��i�؜-���?�v��b����9[�cM ��Ԩ��F���b/O��TS6� �����.;�{0H����GAČ��S����h��e3]���z��RQ�5��Z�"y��5�E���E�2��s*���@FN������U��SHہKvo�,��o�R�$P:�Ն\}PSy�-0�=x���3�hW��_�C�_z'�
UwxU�mt�Hj��"]DI����L�!'�c�G<����xJ\�'.�T+��ڬ��]KK�_�}8�z���<�@�N���^
E�	��J
�������y��_�2sl �B�5�$=�6��j�6�&�,���oyLC��Q��}V+YI8��UL?^G4@���0�0���p='��/�B`\G����{��	�r�@;x�MKpE%I!�E���e�<M?B�`+�/v�&���e�5Jn�����߰{�#3�Ł�~�#�e�!I�Lnʇʮ�Ε�2�5���<�M��x'�������5,:s&��f'������L����þ3���$y��%d���n�P`j���v���fV��%�J�v��g|����@e�PHܠ�V�!s�ޡ�2}&�׳t��
�MY�'�� �U�_:ԏh��)1s��"��mx��Ľ��ʝ-DT�0��}�I������7���y��ޑٰ#��G]HK�����=�� �b:�}i�p�aT�և�����2��2���UL!\pҬ�������ܠ4�DʊXM���B���
�2l�0��t��25�PV?�Ӌ�
S^��8�o��<]�i9
rG����_��"�?s���vB�p�uƴ�J�;MlU��.ǻ_��m ?W��ж[b�2Oal����,L.��OJ�:�����sZ�S�\��������cC�у�齻�:` .A�O�������� 4��P��R�_�!�k�hF�	%" �0cpSϸ*��\,�d{�3v��)�u)4C+�0N�{�>N@&�ev0ȷ�LU�ZM|�A�6탼٦������f@u%]#�Gg�H�J���&4�uE���9�'̇��]ݑ}�f襱�솚_~r�_�1NF^������O��^�'ğ5�624\X�!�����^%���L~&mcǺ�BnP��q��<��Us�mn���-����7��[1�zfF���f�۳��_�|�>��|D¸�r�E���s�&�V�!aN�s��;���(�6��1��Ve���4�`@��I�����u��h7�n��t0w���ry� c=X`p"N�р��:S�C�=�jxN�D��q;Q���""}��4Iȍ�N����d��N�r�:׳k@G�m1譁D���;$��n��������N�{��%x�w5�[gp4n�;��'s�	ܸ{��7~��k�gJbs�\m�k{�dL��U�lFh�BZPc�"R9���g�P�l1s�-�2T��5n�qdӽ�c{����z 'rZ�	C1��u d%UGl�>r�4�?����}��.���G۳�ldQ1�5rB`Ҙ#�{�j�#Ɂd�Ieew�p<�����~@M�QLǪ�t�h�lӸ�ͨ]N��ٯ��*ʘ���l�&�.$�x�<'a�U7��-�֡��"$* �a���f��E�F��u��g����-�w�@8:Y�Vr�ΰ��vhUU�B�Z��'��J{â���^�&;ӳ������j�C7	�Y��Zϩ���|��R&1�Rg5���N;�죩�ۄ�����r�m�^��V��񺤹f��T�>ѷ��4��|��<5og]�O�&��K�0�v����x���	��2��I����*�`�_����YՅ}]�1Nȣ=�2R��㾁.�w��!�4�����\�)�i�}N�q\G��. ��Hhc}'Mc��I�r]pH�NȢ��q�g��5 �c�(!��
��-�wB���!�FAг��(9ht@O^~9b�Y��-mʧ��>�_p���+V��{W�6zC!w�M��R6�<
Oh��.�OH����I����yc�X�4�p�0ǤD-ϧ�
�j'����4�Q-Ű&��R���s��KR���.��9�%z��NY��iU���oQ�a#��q�0��`�O�B���5�Tjn�#�Guӄ�$�$�F�X�|��vE��|�r���aT^HJ������q��$���&�\ǆ��o�&]�5r,�0�2��r��M����S~���_zP
d;YvУ�e��\
��,��q�}:�x3 ���o8\����Ff'�}�~����>T �!��c6��zV�'����[�[N�g�)����s5�s˨�l�2�Q9k�Ȃ_�$��B�"����]"J� �����̳XH�1�IH0���h R�U��!��6��|I��g̤~窩�vǷ��c	�lט"M=�J�ԅ�?'B�ro֤۹cλ�����l��5h�Kޚ��ß�����h�� !o	��_�P%x;��\�Ty��:��U2~x���;�G��T�E��LuNP���do�W��U\(nosE
���d����`����9�*��^ʶ����e
P*����/��L��c��G0+�h�cn�{uh�]��h�?��ߔ
p-�"�VJo3��?�%*�Y?����Nӏ�O�D�rx1�^~���#��L���q�%0��q$r������n����̘�껤Gn)��|�:E��E�{o�酌��Y�𪏌�M��F�?a\Ek�d��F���H~�hJ�)�
\�8��7r'���O���X��bN����a
��m$����U�T���^�T�ܢ���F���F��}�f�55������� �c���"�'o��O� Z������<!��_����q��.1{$��N�cĩ�N1�;�,8J�韀p�|
Uc}vk���D��KƸ���P�#�Ȟda�����0PJ|�W�C�f�KeS)Z6��3Q��U���̖��k��_��
mA���~x�um���ܑA�,^����ۙx���t�`&]�濲�F����,|ЗX�$�=Q��rm���ƥ�ڜ���[��q���P0��ޮ�Z���ۄ8�0��)�>���D<���)��M�>��!�ڡM�q�Nˣ���f}dY��;J�R�9���!�y�Bj�q��=�WT��z�:�7������Cv�ȫe	k��G>̊�B�:�?1����]�Jix��N��x;g��e'Rc€�1�j@`�Pks�X�aXqw��$i#y�}�=n���R�04�CZ(�XV�iH�'�n�$U�v��
6��|�oܓ
�H���f|#'�}f�v
��V+�bn<�-ri�D��_��a+s�9rg�뗠쬣������o�Sa!��X<�� ����Ul�D\S�o�[����?:Hy�AO������'q������,xG`*�Z�����l�>R8C��ߟ���s�x턦�!�C%���mE�}*ڢfF �X�����9����U@}e_ze��7�b ?x�{g&���k����Hl� �Ƌ1�A��A�Y�-�Gg	����&�(�1�蘙��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��R��g�qD�ލ=twމrP���	��� ���V������]�  ��X���-�ـݙ���L[�$۽n��sJ�c�"���ԃ�� �3�_]�!�{=4�y������H�܂�C�y^
�
 ��OW�3�Zavs�,�l���x5�8J�c�1+�[3�<�n�\<f�V_���jiy�~h�L����4�_�%�_��И�u<��d�ޙV�$��2�5ĺ����z�y��`p&���\�ki�f�B�̬Y#�$\y�h��h�F`b����J*�]��v�+���'o��Z6�+a�aI�O�����+C�/�%w
r�Q3Ҋ�3�[�Ƚ�jȠ�D�T�:�o��5�����>�Hk���c=h�;Q�D�쨶l#����R �$����D{':���a5D���:fC�]2���+�(�����R�-~�=�Ķ	�R��1�~�,ͱl�,��G��_�b�U���� ��
����(U�4Q�V=.�a���+4�N��b�/���������_��|8!_X��M�E?J�Ͽ������?�%�5Έ���'oL�k� b��V�n ������?k���}��(*>� ��%��b���<vAݕz�,=�������<�$��O���?dmmam�&Yxa�5߷����5]V��8P�����T�s|�M1B.�H��6��/�Mpj@��.�	a(v����T�#�6��g����׸q��1�s|0�
"*�Ȓx,���ja�%(0F8хn'��q�笺�'wTl��8���,� D�t��2Sx�0 �,H#(m8s+ǻ����qv�d�[�HV�Րj#�|��$�A32�f�jJ8,>O-Ț�ȹ%\�aT������X9�n��5�h�)M�\2gk,����g����n$�v�b�Z��d��^s�tCJ�F:ms˧)���vmY(��]����CK9B��~�T�OH�^r�<F���2�i�\:���摊̾��
�5�[����͆'S��o�PR�Yo�!����	ªv���j�+v�|-k��	Z;�	qެ�-�j
8h�ڇ1�6>�k����$�}��Y�Z���z#���a�}����C���V�.�B�j��QG#����!C0�[�6��ӀL�b�2=��(R�Q�hח�R�^γ����ǧh�]��vG'��w����#��Ι�n�#�9P����T����r�2P��]`��u<`���hz���w�(��汣�� ������o�K��s�^$��ֹQOR�G�i>����@�C>@���.��ݴ��Wc^ڥ��S��rȒ�l��Q�!��X	��(��#b��|��۰�lI>~z͘�E���q��rj��u�]��N7~���c��mƯ���]7Rq�hn����w�R���wz���1~�M�$J�GR5G�p�����ԯ��_��o��a�Dk�f� �ެ&̀u;7m;�"�h��s������mB�ŗ����#��|q�����W�/mG�'�F#d}. rԔ�t�y�Oo��4�w0!`u.%�%�,�*%}ϧM-d���0~�Ƚ�vё�@��~]��Tq��v��j$�wTD��."]����O�
�QV)R���(�c�n�"]�e�ч.l﬘��'��!I6I�[���/N� �!���n&�HL�SD9�h�q��{*aXa�vK��>!t�+���侬���t<��~5�>���dt#9�}aM@�hW����� ��1�u|9V��������|��Pm��bθY��X?��-s)@'�>���οA��S�͛[�H�H���w�4�I�:�t��7��7c*��x�q<-�4fѮ��EA�w���@�녘^M��bʎ�Ay�%�Pg��p��RF�SlY�PwXF�C�#C(�<a�W^a[lPp
5w�8�j�Mخ(3�����Ң��
l��\^���a��Om��h6��Ky:����?Ob����=Ľ[L��vS��u��fe�ܨY�B{\w�W���v���n�t�u64���}d�g��\�.���A��G�s�n�A/�BI������,D͘EH|Ľ����8��\j��E�ā�ڽ{����-��֔0�"�"|?q�KO�ܮG�
8X	^$ܞ���<J��zJ���oy'�Y���ߨ� O�C��[��Rh��2B� �����NV]���6��LF�m�����R:S��`�C�!�(�?���e|�<�B'��t*�pby��κi)��%��o������Π#�M���;T ҦA�c�z ^%��/`�2b8u�!��r��)
|�w.�YY�I�KA2�v��X�;h��q��")8`-4	z!�T�"p���U�OVX�Z�a�sarO���Y���	�y���b.H	2�/�]�V>5��_\Ƚ�f�㭺�$]��|��L�s��{��^����b�G���1|��ڝS��l���{?��3�ʵ+��'ڐtE��c�\��^�xI`6ad�_�����aT�Y����C1����P���àW�*>�����*3�ۻ�*4�����|JZ ;�����K.����\��^�A�^��3�4ċ|�%X9���Փ���B�$�saY���m7��`���;�G�F){F���x P���}rGu�S���PT��xt��0rj�����dO�&��|+z27?�ݬ��0��zM1cV���~|�2�� �%��Ou�V2����Ĭ�㈲k��b>=e��v7�������A#iПY�ɼ�YMR����[�ڼ첲R;�PۋeW
[A�!'��L����I�T���2c㪲�S3���2h��0��TÎy�{\p�����Y��w�45ufy#����t7�ph�Y)���\�ZB�]�6O�����H����kgw��	7�&3<�Bf@U���s%MJH��n'K�	&���Q�t5��Da�#B�9�Z`���>��$3��و!��­��f��o��"ܺY�6�Gۣ{�%��>�k�7����q[��9��c^���(/Tm��4B_�#݃@�e��������Y�W);�yX@ښ�2i���b��gN����Ѵb$����@����M�X���X��Vᬙy�y���Y�E��q�,F@��|]�ϊ�����
?S�N�_��zȎ���=�G��(�Rm��������r@x�9��ݳ�^F�I�Ԣ�9O2Иa�y�q����r��R����(���B���]U�M��n2}�},lf,f�� ��>v�{Z�׺~o","T��H��N��-��(q���p�ͧh�nnw��I�d���&{�Z�Ε��zb���I�6>F����Kq^�2�Su౬o�. �R�8���z�v%��pk:�;y����fT����FIeȢ��,x6v5�h�m��3i(J�a5
�4��M���dB��s�Ƒ߃�:�NQ�淂�>�d�}��?Wok��M����`V:q�k�6��}?�_���di��s�Ģc�V3q��J���s�-m�i�^������8] ���<ɧ�ϳY��L�p�s��L�u��{m<����k��Ǌf��؉p���8�,7oE1G��$�1��?�F��M �4밙P��%��$�O쌀͘�{!�d��Mɽ\
��,`���L�綞Bؽګg9��c
̒�X��������
dɹ+&j������F{�@����3N��ƹv]G��\�*u��z$02,K�Ys�f'��v=ߛW�.� �� �_�5?T�+�D�xq�;�]<m����4�/��0y���+�=�m��H�r�WE��1�E[�h"�9��'�8�-�I;ob�E���U��ܘ=�sY��Z����N��"Yt[�Iøz���v�Ό���w �
�\(�8���)l2�V��?���;��O5Iqw�(N�k��!�	��P������-;+���w�x)��=���I�_3�?e*�|:n�ԛU��nw��K)�[����F�-���{��L�1�7pH�����!�n�>4����Xv���̒d�Z[D�ߞ�Ľ_"��|�6)�-Gy ^�
���0�����V�k~�pߣ��"��>��|]Na��v�/�������a��'x�T��H�e����F'~x��#< >o��}y�ݯ)�W"N���7���hEe�k���3���nZ�yޓEd��7�㹄?%�����|[M�%�
���	��e ��4�F)�2"���[�`H$��O ����l,<ע�z�M)��rv?�hM
��A��솸=�g�(�d~�F����K�Xm�����k���L�ϫ�`�j��lQ�ź��B��s�a?�-q�Nڻ�i[���c���O�E�V/)h����ʄ��r;���¼�o��O"�)Af~&��ty�.V��@��	�4��X��!����.���Fkr�G��i��y���6��ϩ�4f�Z��s�Rv��M�/����ɱ\�[g����|\��옽?�B�v<X�rι?�jٽz�{�X	G0é��z�h��5k�,��O�C���Y'Lb��q�Z[���t��ǳ�rgor%�}K�*y$fS����H�-[�{<�\\}�5츁V9Ǽ���:o��/��y�Ni��FE��^��R������C�����O��i��i�� 7?�_Z(�h�&3	��=��j�@�OΦ���ss&̡�y>�ǳ߹��e׷���^��#H��a�*��@���v�����������{t�r�O�׋�~��_��/�K���E,�(���O�ǰ2�+!z��{�܂޾^ #��w����?�w앧�)����)Oٞ߸�e1Nûk��8$fPO��W�>���v��qN#������A�W:�R��ɷ,�����u*�E#�@-oG����j��͜e��*�zaȫ]D�G��3�N�:j�j���r �%l/ʖO�#�}�)Rj){�:�#�6���vϏ��4cu���_Y�F�5��>����W?9[���Mu��9�Z�+��w0zԞ[��I�y�˘x�)��&�/+��'�%��|��Z���Fܱ�Hѕ����;l�?Ԫ3>	"	,�Y%�����M����a�D'�M:�=V�ĸ�����A�	�ִ��ܗQ��6���z�����OJA�Y�C�8E�P�(�W�5ڤ�I�7D��k�����@���Q��aB&y:����ĄC�l��
��r��E<M+O%0�w�/�#�F���\n�X�,�.W<��G�����|� �z�ad_%ь�8�#bܢُ��q=58���5%�+���sZC�Jr]�<�xlj	���_җ��L���~���]�t��	r�ܳ���6�z������(���5)ve躥�!)%��?���W0�%��7Ӕe�+��q�1Z����p(K`�/���a�α�����o4�l��G���7�5�rGy��<�b#��g��P���С�Y�w�+��A���Y�ǐ���������5�V�v�\�s�93�X�l:�(�*���{���Ĭ
\]؋�����>�����H���[o)�&��2|A:���׍�/�D�@��iցL)P�*t����;�m�.vh]M?id\.H!��!��]���h3�v|B��a��9�0��e�l���5�m��B����R@��E���Fd�K��-��kU�8Qn��N����`?8֍���'�[�G�͒<���N��vf�p��$�3jK^'U��O�4�����~�|o=�u�մa40rځ�U��s[�I� �K˪���:��[J�r<�Ak��G~���%�u�jF�$��3�1S3���{y`lwjW6����B)�b�a���Ev��i�K9m��[,q��hl���C��9t��'��k��y7���0_$��|gt������L���@�8��*,+�ݘi��y��Jr��E����u������ q�J��O������O�a������9�^��qbږ��C���&�U�}�c�����ψT�����A��ԙ��,��G�9n������3��s��Դ���7jʐE�{�
\,��v�y`����	݇�w�$\ss{��r~M�WF`�Y����Y�I��&}��i���;]w���G��|��Q� ���] @{鰧g�.�ʼj��	�l�.������ e��Td$��~�&l�+�*����
�� ��,�~aI��ʼ�5��������
�%`��I>}c�"�z�	�n9����)�[��Qv�e�
�Y�&_.��Y�AQ��Jl#bH���ٖ19��L�*;t�j�
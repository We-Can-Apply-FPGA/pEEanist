��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gs��.?7z�}�����)��T}k��[o�E�,�a�w�v��6i^3}��UqJ��D0˫���X5u^Ժ5A��J�����q��H�q�S�奈��s냠QT��� ��&�,�^C$0�>h��9�O���G�$���Ր-�a����7A���4���-,�C$��`�h�!�%�k�Y�A)v�s�'�0b�K�f�i�z`����7��6]e�����Lx��4� ����nu��<iL˼�*�et-�P�0�"u2���V��_Tq�*��V��'ߟV�[^)p���x�^@��J��.���]�!����Lѩ�1�a8�xM�EB݈~��'�'-i�����t�K~~p8nF8{$)�|�Am����[q�+o_�f���9������d.��'�@w�z3��K�{�LWį�鼙��W�ܯ��=5l�9�Q�6c�����ai�3�?/ޗ�'���}}kK��K�n_A�.7���M!M���9��"�t��K&���Z\�z��(�<g��l�p���>�Q�A���Q��22��+K����6���	��й���������\}����k��HLz�o�Ds��&���gQ�2�5�g��{�
�!+�`�#�� �2���^�c��wk9��������	v<�W�eԤ��*��a0�K/2Fd�ƶ��S���r�j����������N����\j5��1I�(|>�M�0ʿ���,'A� �>��R�
=��2j�0��z}�qYK�\B��Z�\
�Zآ�(��)Cn;#�"�3i�KRe��CB�X��V3%˕`Y:�>�|g`<�[�Q)	dSP����Ģ:I�����^���T�7���7��ug@V\�v��2�a��JQ���o��bS �$s�_�H�?��ei����)��{Cg,cpоn,X��H�z\��T����!�������)7��	V0�,�ƶ���5��@���W᝱�}�8�N�u;_W��Uv(8���[���I\(���܌"Qj#�N2�n\�g��j��0�|;�8�N�[.�ה5V"�޲o�J=�S���9h����q~��[.��Og�t�`�S��O��fa��ʲĻ���s�:��7�N�j�QW�����-�2����XY��h�ʕK/�|z2�"��A��5�d�b���c��:U�U=R#��[�I�^�+�߳i�k�e]��KI^;�̊�r������y6yO)ά����X�wi��!��'�鄗�%C�mT��СM�'����m�Kr�0�6�vP8�N�[���uG�㧞>�&�R�)��yW�)�8�G�֚@)=��N�w�X��7�'�Q�P�"�?%*J�1m�&� ����t4�|%/:�U�MI��tO�&�,��h��<�g�<Q����:O�7:2��^zf�ɕ���-��b|O��;�w��x���T?�ٳ1�lω����[ðɘ{q�����^��ɀU�G^�F���C*�*E�O�l�\Ғ`d���Z�J�
�����8C�۽�G�΋౧Һ��~,֙���䨫�'g��"�+�h,���ǚ�!�tߎ�ZŗW㗤���B��'���hX��
�(-�x�f��~�}�`�BRixyx�K���j.�#ҵ�h�Cl���q¥�����_@ncz���q<y�A�J�g����v ��# ^���~��v�,��-!⮩x���iS#���s��̱(q�$tˆ&1]�.J9�L�6(9�X�K1긃�+�Z�̱�s����=�]�,��q��k��,�D��-���xJj0P$�֮n7��2�w�<Y"�h؆��mO0����6�*��?ĵz�i*:��JGh8�?�F�:N9�*Ns�Ⲛ���?��}6�>�-2.���s��XE�-ig�E�	{{� #v�ѱ��VlS��AigY3{��A�,9��[;��w�M�^�	�| 3R��jl�/6���D��$��as���t�%�)J�����e#
i�	�ߗ3�?���Q*-1�(-=r�y��Ȟ��q tS4{��z��N�,!�e�hħ�\�,`M�P\�A�>/;��ņJ���Ǔ��K�[:Z(�LcKpp�>J��vb:�㼖� ŴE���^IRN	����py�t�6�$�.��=�����aQε�<,��#���x����}.�2��:��\3�j;y�[��$�R�أT��pΕǿX1`v4�)m���v�E�k:����dJnF%W�W��hM%h�`��5͈݅n�^|�H�b��L��ZLR��BuK_[�rt�3Y{j7Jv�Z/޳�*�Lx��KE��%��w��{�� $�wm�V�ޣC��� Z&7�_k�Q���f�f�]��>���V�t�=��Ĭ��_�a�,�@�d�0�� oD8#w�<�Y�����)&�D�:n<l��o�N2@U-6��\��O�[���a&t�C�4�T�8&�6�t��:rN�����>�\��I����Skl!��lE�I�;.X�T�Ǆ�d#lJ|�ase �v񙤾�V�HLNʎ<�����㽹G'���
l0���(����C�H�fPT1���5x\�a�i����8��F&�������樍�GZG�ж��Rgkc�N��+H9�͈ܥ�D����7���"ᛛ)��%�pP���.�ty��Hy8���%�7)#8m�_�C����=����7C0����b�)�ڨ�r��Rۀv���
�l2�4Fh�ZUP��J	�)2p2��r�ˀ���
�
�������%<"�J�R�!s��a�-���D��O��M[뼇Zn/DX;�r6R�:i��~T��\?F��|W��?I#P�3�r���l�[\��s�H+t�ӊ��q��ޟ�K�Egm�_��_�,��g��CRRc>�����o#��AL�� 4`���)�6R��{7�>����'�~"�DV2[��wN:��2��=�s�Pr�+�%�2� ���rdLU��VoWVx���Q�%K��Ћ��``ş��*��HZ�C�qc�������'�$c!lX���N�4-ND��[yE�-������< 
����ya��,w-�������s�s/�gc��3vG������!25��x��͢@~����&������+Ž�U`ʃ�"�E�g�M�������Xm�z����]�#)\@E���p>�X��W9��n���	e�5�'W�r��p���lnɛ��ϓ����e0�s"���(4|�[T���E��/������o�S�A6V�2�d�Lw�]�
�:�B�]~(T�>UX{�P���!`V  ��=�����}��*��G�A9��T�̧��٩I���`�nfv��}��g�����GL��=�׬�K�z%R��1���%�C�L(P��\�tW�=N�]ǔ�f��. S��"��w����q��%�OYB�f�7�]dz�Kl�l�X{
�D`?Bd�[��dpc��i�.�6z�t��r�J\wѰ���k�nG(�w�e�	�#�5�o9�
��m�T,��r�$L�N�'�y �����n�iӣ�f3s���M��#���P���#������SM��)'/�u�vG$�)\���-{e)�玫�(0��	��6+"h��E�f��Y����j3�<s!�NN�>�3���Jeo�"�X�Q�Ez�ps��?�@�z�z������V�>�s�+(a7�J��"���"�n�^{��l��D�S�����Ԕ�l�z]�:�ͽG�_﵌L���=G7T���/��$}�s��~���#Aq�!���j�c�!���u�y$'3�)��模��[Kq�9ׂ�G��pr��1��
�J_2�!��+T@�sv�U�d��x��Z������}QsXG��s�\^���B]4�;Άb�fB��e��� �q�����Z5�=��5��Y7�����D�e�u��.d��D}�m)��|B�gYW��w6���]-���'�V7Zn�
���O�i��6�rŒ�֘�3�l��3T��p2�
�����E�QL\�P�V�hb��
#��frsZ{����S�ƅjT8 ?��Z��R�݄�Σq��Ny� �ИqX���Y�<p׻@�R>��+�3�%h��i�)���A#C�H�>�̣�jG$&���r�����սP,�Ӻ�I������t�d����~�@�-�!u ��=��}ޥ��9{+�����S�ۢ����W䇹�S��)�P����WXa���|�r��]OǱu�<]n���}���D����͜&}kyK?��������s�U���Y��C��9���ի�hYGI80rB���VR�����P�����ޜ<���l��w������f.;��3�4+��sl�s�`�0�l�h\7H
���������[?���!��҉��(����.��RL�rr'F뭯*��D�P���=@�oyN~��GՁ��k?�;��5��9�
�D��W��2��kL���V9���_�u��Uܨ��~�x^c!�X�0�>����i+��7�dm-�ɦ,�����[(��5q� �":;{S��D�]����y�'.��O��ɘ}'��,T�%���[H�i6��|ו�V�G�@#��6��	��l����d��Oy�[�1l�xn� �>�=��"�
��qѬBh�lR�|<C�6^?��6�9-�"o].��)�"��� .H��2�P�3r��_m��(\����<���]F�Br��+~V',��:Z
=:���;�~F������g����V��1	@����8%�n�@vc�!�}�w1����E�7�B�b�|ra������ �;���ѭu�L��j��$Ρ�?iD{z~\�|�=Z�)��am$=�����Ά4�e�]���*Í��b�U��G俒��3���@<���
x�j�1�!�7i�Q���������O�"L�k�&g9��	��	��bgp����s���T�6��l}�$%|�Ϥ��	o����� J�{a�@������,���,�(f��c�ҥ�)����.N�0$�=��a��7I�?�{�����U�U�Z9�JV��S2�������O&a�9�p>�e*a�<��
��'�����B��\S�kD����7/<Jˆ�R�K]����|��V(�`7ZL%��qJ�������[�
�cin'�dN��^}�yJ>��~�6wz��l t�ͤR5�{��1?����b'�IV3�~}����QiQ�"�JV�=+zl<s�H��m8��C$=n�G��ZbE�%wx��|���+t�8x�����z�*+���I,��◶-�c��ؼ�K�Pj��2h��n��<^��"�c~�Eh���b�d�i���6{I��6�
�F����50�F0���H2mP?WVK�����7J�������� `g�q��O��U�2�(�% <\5E9��5'�Qk����\�=����^�-�;�I�ަ�]Oڂ�z_߅���ӽ76�lS��3v(PzE�n������"�%�/Qs,y���x-��I^�Vh����9[��5{�WdqS���ޠ�;3e�˟�o�6��[&zO��D4�;�0Mx.,�=��*h$��-�[��� �U��������ڃ/h�B,:
�����]i��`݆��pV�h���ZB|^��q�EP�~)���6��������U���&����[fsX4� ��Ev�%/p�=�> N𚲸{gYnD��5����6b6"߻rKs��.eF�Z͕GL�#��L֌}���� E��������`�hx��!4#�7�����ٌ�|	�&���N�-?�x�V3bŶ�jЍ���pO����zȤ�<"LV[hZ4��wP��rfT��BC(�{���I�#c�6ƱpǁB���2��퓡����'����^ �6ХM)g\�%B�sG��#�Z�Wg�a�l�l���OO�R4�-����Ńx��\��^�
6\Pf���eˇ���}�V��,�eJL��z�L��ޗV�:˟~:�n�2�W	�y�4㲍���H��`j�`[W�?2+5���Ϟ8�M݉�kxՏR�J��ݪ5����ﮞ�XjZ�i��EbD���Cs-�c�x�����T6!�����/�;�m��E�t�M�M���,�����FW�Cm!��H�+2OW��;� ���$y��\69N_�Ň`qѷJ~�[���<<���*��q�H��cb��YTk����
3R���K/G���q�C1T �M_����lCA,a������nj	�_P���>��c����Nݣc�a�����C�I�ЧjG'r+���ד������VXu[���`2:�������,�^���<��v���ش#�Z�Ʉј�����J��3.(1j����/�l�YԨ�0W��h��?^Dz���rz�1�5�`p� ��NЖ�R��4��cM<vW���h@�6Ǟu}�f�i����U�p�w�q��5��U��O�)�=��ۃ{��d���]�@_��o9D�i��@�rS<�}��6&7����- ���E�}f���5@x�CLI��c`�F�߶�]F��aW��%� S����n�>:�g���s�z�&�6��yg�s[��'֋�˵��$w��/�3S��Ѕ�uݕ��*�Cb���%J�O+O 3D��ON׊���4?`��1PUI���Z�WM��E��[�dZ5|A� \+�+f��������^_�"E�0�[�Xڑ���� �E��fuk�Lk�!S&�55��7�7���_�L����k}��]5H2ᡢ��p���8�{���R=<�X�fԳ��du{?L���t��B����8�?�:����b��?A	�ka�-p�ew���b�l�Q�\V���7�r���B��Tv�F	���uW��R��b�P�E��Dl�߼��#d�9Z��G:W5�\zɶ�6µ���N5���=s����e��O|.���zp�^�K-��Ʃxv� ���xc��/�%_8��i�R�:� �N��rR~��HI�R萁}j�=��gu S��k��!1F�e \��YC(f*!s�+y�Qt"N$��R1@*$�ڞ��<�@�;w��4���3�+���38��%e�8���3�-�ݏwʪ`w\2�p`rJPL�tf�9�7ĤO
#o�)��3��P��U�d6���Ly�5�h�����!�:��V)�ks���U�L����g�o/�� \ ���6��1Y2ث�4�!��r�m���ە��~3`@��vulXe���`�J�ف6��6rG[i���9y�DQ�)̑o��G)�%^��Vw.�k���tF&��� �	����#Ln���qV�$Nq���8����&�o�-j��4 �1D}��`2'�'j��7~a��C��y��Ӹ@��$i�hQ~bdi�B����iP޺|�ު��A�'lD�y� E��h�����PR����>��c畊�����d�*D�xL_ë��˟>F�,���9�]��Ҕ��7{����W�0a�gI�-�����k6j�����nF���g�������y[�c���~��>���:�)4�7ک섲�;@9�=~S���,��7d��*(]]#��J�d�6��Uv1�ĝ\�gF�9o, ^�v�p�O��$8`8�+h*N+�#�f6_%;�����W?'k"��H�j�ˈ�����]R���2r�>�/�s���D�0J?}�m}+v~�=rо^����ߟc���!2Dx�j5$�M'3��
��G�rCWꜘ�/|���i��<\"���+I}+ƴ�#�MÂ�gm��(�z;f��0"j*���0<8C���r����@m'ԡ/�	��|ئ�������?z�oGȧT��\߿JR)�Ej�ϓ�'��~�P Z2�ҫ���g[�����bX�9Ry��*C�7�rN^.6������v��e�~2�0�>\�l�Fc�a��`���A̣���D����1��4i�
��vAP�,̑
ԋ�^�{��b0uO'���w0=$��t�����*oљ}%�t�M������e�t��#i��jzyZ�̳\�0RƹM�R���u�,��H:��D�h�Ti���S\�l���~F�
���#�&>m�R�����*��^�?���A�����k���=���,TiA 7�����糏P&it���;@�S-�V��s�{�a����[ȉ���P;�{CI���%�h?"�粄��Τ�J�~�2��l�ªE��xP� z���C�\�V4B)����F��#7�'�����22��u(ݟ]�Ɋ�V5��GES\��i��IE�1�����}d�����c��ۣ���, .�ng�j�Z��X��"�;Q�[�����Zj����L�6�>�@��..���V
��d�`�V�y�h��QjK!�Ϥ�d��}�4�������#0��^�	����C;���ɒ����z��{0�R���M0�>���%��ve����z$���� ���(����`�B�r)/5�G�����#��Zr'i�?�rѯ*��d�\DK)�\�m�9������$O�&R�;H�ԣ��M�qR�0�)Y�mx�����%��#9�pA�5�Qʋ���lD�X�
&�Ɖ4u`m�L�~�C�Ad�@B=�*FQ��cW���y�P�%�uD��<qT���܍�f1���@U�*I��5��%H� �j���Q���V�)�=w���6��Q@~��˻�R�!m�%E,Y?����n��z#��J`���M��L��[&�(D8��@:�F����y��Xv8,TSz�
��Q����}��b�m/�L�4gN�;�o���o��?x��2_O���WP��Y�y_��s���:� 5���`�T�A�Q;���^8�O�LE�����,R��`����� ����Mb�)Of ˀ�r%��5*=w{W�<���"�m�7I&9�P1����4Fr�?�\Y߼�^��!��/5�w��s�:�F�3�|�`��
�@����JN�V�H������
cM�(W����a�No�df^^W�G��"��E ����4����3�,�b��yN'����
�F�M�̰��Zq1������)�8���Z�F�i��߇d"'��[|l�lx: Sd��������h�r����@�0e���uB��7ئhb�UY� @βupĀ`9�@��ɞ��x	8�����S�-O��$��* ����?��!��hVX{���&!h�������n�=z�m�8vs���Т�י�s|�h����٪��x2�/�L���\�U]�\q;��f;�WHo�y�v��*�c���y�	����U�A唎��>�J_���b;u���(!%g<a �$Yle�q� *�{��G58'gj�H8�.'�c'�l6ʁ�dPn8~��o�麹p���|rͧ|�&݀�l�����[t�QoC��Q�'���2�k��J���͖�)�\v�b���ʈ��=b,(\ �l��r��?'�'���JS���h#�cX�z�J���G�^>��������y��g=Z�]A<{�+�`��<1��"�Z��'��X�KqW��S�h��8o��.1rD���#�i-Eߝe�B������K�sM��ݜ�]��ْn�f }a��3h~��K? �����v�����F����T�c�"^��	u���
0��̷X�,��f�S�8E�����	q����ג�G	�����R�-��k���j��N�f�5�l���7Av�Q��B�c�o�l�����Ńʇ��͝�/���il��
��?b��*]#�ԡ�j�U[���6.�}�w�s�]�vy�^J�ճhNU]�0Ͳ���R�Č�c���/������ۈ�i���-�25A�-��#ϧ,k9�ua��;�~�x��m��e�*������G�	�|@8���z����"�Wyi��˖����>"%���p���ҿ���|�"#k�p8�X;�y9w�"E�"�j�ߟmfzQ�C�0�1�q�N�� ��]���J��s���H�k:�t�j�����Pc�c(t���D{u=,ҁ�[82!+F�{�!U�~E��v�]��"'~~�Kxq�� �����G2��r0w4:Ö� �v
~Ѵ�7�T���b�'8h��M`���[��?�=��;�4\n�|���ŠT�7��H�����q�;�����~��3�҈p��9���'��`1?:Cu�@�Yķ4{��� 1�H��&�g����++d_
�8�A<����=�2n�]��Z@�*K�����H+�cao��<U$r\��>1�/�����L��Ct�-�z����_r�$�R�d�����M)�}�1����7�*��'�y�v:���@��ٞ��,��Z^ɞ� ;>�L�â�y6��3!�L�DI�	x�$�9&����N�MY��md��n�ĘJ
L�_��&�R���ܯ
�����t�>�
K�n��V�Yv+�1K9��� ��u
O�~IITD����j9n.e-8��t��E�4�h��+7��#�/ s�$7�r� ��4����N$�AY�a%lv�Fq�]��	j56�썰�8�h ��\ӓ��8009��t\FA"e~wڂ?aTr��D���nXv��.��{�%���PU��p��u��y\�d�F?h�Ɂ���?i`jXN�hT�i�n�y~�z>C��~K�1l�T�W5��&��i$ՠvsn%2��<��m��U$��n�������&WP��L��ۏ��l	���7̮��7{<N.H��o��[��0��#5r��e]<m9���H$�*�h#��3��2YL�t+Z���2E����D���X�ȫ�����N����H��a`���J�m�������֫�lP�8�ρX�3�&�����Pc��L����0�X�(�,EU?���݃�wF_���3�S�����oP�r��3Wԧ�3㞠z�LcyF�[ɓ�⟯4e;���pAj������
�V�vP�x����Ÿ�tx����&��l^�ޅ�m.���9����OV���q��Y6�3^]�F�	
�^g��C���'H3m�kc��D��p��cdt�ȿӻ�P�YLA�\����rGUW%	��$��L��yf.'N�8�A\|]t+��DC8���3�Qn:v;��K�����ﵿ��T|�^�<_��Q�ݙղ��,����y�%�_�5�����]�.*/By���f��U16��=�tgl6�w�D���Ѓ&�<뇚��L����)w&�%��Ҿ�3Q�65���y9�-�B�+����KRƞ<�(WU�E9	_R4݉�J�b�w���^Z�mZG�*ɶI̴cw��A��B���J�=��I�����0�`�ڸ��T�
{�w��x�t}��O��/W�%>2�������77R��Qb���|~��~���b��;;��YX�MLgw�&n~fA�#�3��7:x�h�s��"m�Aƍ���`Ld��sd�C/K�'��1oǇ6��,K�����R¦ʄ7:��y�Ḽ�'�#�z$�q��l�\����m*����D�y�{۠�քB�P����*�4�*>�I�O�����f߄4�d�*�Fvq'�~@�H��]�V&A�����;��ު�j<�o*���u���Gڶ�j�x�7(��n~�GD���o/�v�_W����B����_��ad�:YV`rH���,l��L��z��S��(j\�763]5����G��-=4	����}#�C��_hU����<q0��>.<�#�l��-3�i���z�jӊ���֞y���a��<|d�d8�Gw�m.��t���'o��(�b�����U�L�CQ��iA��A'dT"~�JhLTn%�I۰
6�4��)�J�J*���~����꭬���;y�(J�3v���t�?o�,���Y�*#�Ȥ���s��T`_��
t���ke���/���fx_�.ٿ.Rp@�(¥		B�D\vA0�h֤���yv�
;f��~=lC��A�3B���p`�"�v叹S��f��&Y�bnc�D�	� ?m�վ���.G{�-s�-&�F�V0�Xף�����q2NU�D���,�*�Jk���l��`�E*�{B� �#�'��Z}���U/�+���A ���^F@�ݘ��|���n� ��?��D#�T$R�М�ʵ�u1 �l-y�T��e@�%�;��W=��^��~bƴ�;�_$��u$Z_`8u��{h�J��A3�]�Y�O�i@?�i��Ȭ�ꭒ��j�$����;ò(?hZ�4�;��ȶhdQ�l�3��G�-6�y��`Uŕ�([=��~�����i�ˑ��D�6v�)Q~�;Y*���^b'���BZB �@��"G�I��L�V��4��L�Y�z�I��?��L0�@?��2���2<;�&__�;nQl��#�a������!=�N>K%��9��YV�:gQv�����E����a�p��P�H�2C���;���Θ ����;Uh%#m�סì`��Ir�ޠz&�M������Y��N�j{P-�E�N�Y�
wf��-x=�T2{���i���0`?�Ek������\HE�����x,g;\�ɖ�������!�(���b���	c�nȤ�4���ڀu��V�D��0Ü�9���V&P���~!U��HX��
nZ$�Y�/y��p��/��>���_��!�bF�hP%U�D�o	+6ٹ�Ko�:vK�����uY�6��.ڴe�yj��Q�f9�M��&ܗ��2���)J١��>�&`��j��A�?�aH�Q�$&�����Dޓ>���������	�6evk���x\�7��:P�,�1U����`4$3Iȭh6�^���
�=1R=���s-G3��u�@맺\��E�[�G9-
htk���+���W�i�Y-�� �R���6���lP|�u�왭6��1X\�-{){����o���[C(�Sŉ���V��in����n���Ÿ����;Ӳ�Xa�p���O�)�8�(q��	B�tC�=��8�}�ר�^�@�AD�^��覽�$5ug�5����,�n�
�T^g�^���WA�ph�{�X��y���q]?d!�Be����|I�v�2��Z�	�p��ܻd`������0��m���g��`���*�(�+�3/�F�==�	j�˪��Q�8�/�����jaG2�O٣�^�J�aW{����42�Bp���{{@�,ךY�c�o6�z�7����p_uV���gN�	�7�����l���>C"�+2U�P��	,���ntTʬyY� w�@(���e�3E����@}����6�nH�YC�]Ժ��E�*��
���ڒ�*���L�V�/��h�c�K��f^��[K�z�IͻJ5��c�/��X���/y-I����w�YA��=�*b��IAv��m!���3��fǊ��	�(��dx����߁�Q9p���B�Q���ٷp��?���Srr�J�z�<�yRr
����P��tΆ�ܶ	�A�CΖ
�|�Ǵ[ �!��&r1�ρf���M�]= 	�!���&�k�1Q X� K����|Ek�!.������N�}x�A.����t�fl��>�����������D��!oRyn�<~ɰ���w�ev7|P��ui�"��������2f�N4[������IgE�Ѥ���Ǳ��f�ْ�RJ���>Y�ч�&�<x;�y v'C26���}�@�c�tG�l�bU)A���#ڵ�
6�@�*�Qs�μįc�fl�]EW3�r4kX��f��-l�c��S}����R�b����؉K����!F��WN
=�A�׀�>@ ��n�Vj���A*�t�\V�<i*cĎ��>#4@c���b��3�V��ǬvH�̚B�sA��xn�=+�g�v�T�9\��`vi	��r�v���#aФSȁ�hZ�?כ^؄"��$T;���^���a�wA�N��S?g"��I9�˚7 k��6u�5EK�s�Dc(8[	�_0�U�X����#�8��%�U.e�k.�$�,�G�B��h�(�ݑXA-z�F��p�+�\�6�nЉ�A�v1�]TW:&f	�����8�`�Q�N��6s �uz!�.�yB��z��t-M�ڻ��x��|ڶ�|	�"Pq���'���a꼺��ׄ���5�f�"[���Hr���R����U_�F����q�E��B���r�E�6���ӗ7|�a���l���2QE�qv�~.�=<��g�%���
�z�ėH/�5\�_*���i}�������"�/AVǦa�O>�m �*��T��e��'�6T��.(i�=J���5��x5��H���(�f���V�:,��R'ѣ-޽�A�\m/�x+��C�S��^��d��-�}c���/_Z!ٗ#���ލ���K����$ z�"&-���������|Yb��G������%0���>��~a6�D�A�NN�q}a�DS��ND�vb/��rl%��:Rq�^R	�RRy���#�)��!C��o���~��%>��c|������u̷��}���A[&6��S8'�8+x�DP�Q�cw�_�����w�����K�k�l�{��*�A��ͺ= ����Vċ"�੒�F#=*����5$�hUj�N_s��d�ʢ*���ׂ~$]��-��53���n��g�P��9�iX_�<���S,)��VD�eK�0�F�d�փ������2\2��9uU�
��)'c��ݍ�v0���?������� ���!AM�
^�����#5�,b�������'>c&��`�{��Q3�R09<Q�f5>)���[S"+i��N���D�Ȟ���Ǹ��*�����'F��=�MH�W�r��3L6�ς���aD��������i�~�R�l�9+s��W�(�PX n5�<������Xq�ǕhZ�'���Xu40����O컇8�]X�e�����ϙۖ�U=AV��5l��F/�/n���oG�z���2�D	�Z�|�۱�c-�Q����;�\���_vu����GYAY��^�Je�*�m"ʡ�+�U�M|��{7����o��$�{f�8�/�&���MRH����ñ�mQc�����F7���@V�^�I�>�E�~���2YDFp�����drB��RM4����di�D3�]H3����6`�:����O9�m{=��F\q�� ��K�`���ShJ��>��v�[b&�vQ 4{�nR	~�E�84c`�Ώm��z>���h��ꆻ��$��B[�m��V���m5#��El?�Z����-~L�_A>������'c���%(�7c�/�ND[.;���8"��r�*(�G_�UJ�lI.��~�����I�5o:u �Sˁ V�"C8V`����������w�G����
��r���PO��5��I
;"�ٚ �^�,���ȒxN�U��$�6��9S�r�0��H�
s�G�Q���$���I�
��������I�bŝ׌��J*Y�;W'&�r��I�	r�F��h�P�9�:W�{�Zq�9V�ǔ,Fu<V����g|ؒ҃����`��{�L����T��-�¸��J�֢��a�����R5�����mB\�R��|�w����H�`�+����az����sB�ӵ�eit� ?��^�ܠ�j�h9r�ɿ~Rm�yf2P�x;Kgz����1u6��$Tğ�����SL5�Ӽ��᝖f�~i��剩�l�yb5K�Qޣ޹�1tHO�]��n)�6"���l
$��u"�	������-��o�<��Y�G{��Y��G�0�2�,6J�~,KF�s�xG��|��Q�n�C��?hj��w(J�-�/VV�z&R�;�U�˩�}��@!�IR���{�������*�"źe1�l���N[龛��� �I�*�P�ם�t��ې��'-�F����5G�Jc�wD�-7�Lͭu���8�A?s��!$8�8C�N�� ����XʿO�s�[�������2��2H#�Q]�pu՝����j�~Fv��:9����!�ǹnx\�����M~�8�;�Lo��O@'��������MK�͆���ԍ?�'~lX�Lh٨������� ����r���`tKwu�]v0@1K���e�}��9��e决_����(��5��z��%���wOТg*N�E�W��n>��-l9U
��>GM�}�lf{�

��H�51ڣ p�r��O?��o5�׿�)��i$�47�6�������b1ڰ��F�iiz��Vng	@����e�=��f%��G�<�<μ��������!N�t%K	z5]�]��~��㏎V�Z���r
���2g&s� ��=����'\�O�����`�A�F��k$�>K�]5��:������&"���T\o�����1I��i2���7��)��� in�y�+R@hj~�u1o����l�Z/h�h�i��'�W`|Z2 o�
t�;x�}�2�{|��v��WZ�dgѧ/-)�p�&|����J�X1bIׂ����H2:���O��u�Ċ����̩�`��C7Q�c0�l��w��[�C��+�Uk�lSa>��3/U� ���pX���d�郡�Aha
EC�u��o)� t�։vf�s��V7&��Q���W��熟�ݒ*���
��M�Yxʅf��A�_i(���ÜZ��[���bq�Au5`p6KG��d{�&�K�W�My���#�Oѻ3���g�a��zX��v��8k{44�"CTן ����*b��;��+hy��`����`�^�{�G��e�eo^�@뇘��(U���يq-�4~��(8��U�b��s-�9��U\�Dc�ߡB�,p;]���I�_�����}�=���+\g�Z�_t�X$T>�8�����J�/#��ڷ�zֱ_�n}�����z�� ��S��Ny�Ko�1�A������c�nPL��ۄ����Y�h9�v)��)�b���"�Ȯ��{�~n���Je1Qc�o�r�,�܋��D �����(\��<l�&���
����1������bgo3O��8��?�Q�g8��� �0�b� ��x7c��a;�/,��}e̩���`|�0���)�r�[[T.B�Gf��BKO���o�fA ���A�f�#Z��7z�-� �Ŝdf�Cc61��k���ųBՎ�";�/�w����ZZ]�yl���?�,��RQ�R��ü�!�8�_g̾�����A��!:�,��t Gw�T�������Ԛ�#h�H��҂Q�Gp�?*w	Y!��Lṳi
�=�����]��,v�9�C�ӝ�`��̩�RM�ݛ�8r�,ٴd�DI�{͟�~
������0R,��Zz���A�æ��b������Ҝ��ı��S�yhY:�w����'��k�WR������P��f�u�ؓ$'�-K�o�t4{�]<XSi�@Ȃ_���]^_��'d��z7r*J�)��U[������y6`�z�S��©FuH�Z��&{mai�4�˺�����{��U�N޺;��mev�@��y�{��Զ1�Z��Q$��n��H�d@u��p;�e��xk���������GIY�eN��'a'[
uzP�DH�X�m%2���~�yF�����a��㨽�C����u����_>����Y�%��9����Ȯl�`"hkz���F+-b��r�Ⓣ�0?��������͋�ڞ&=ٲ$�A���4�:=��sC��y��Ub��/� Q�w�BTXA�S:Ծ��>ft���m݄b6�Й]�<��$�y�'�%@M��d�9�>����>����sz�<:ɚ�b���"l��@tB8� g����$J�@	�&�@��"���3���b��3�W�]�C1XsF���jG���|gU
��y�$>���3�w�>h��>�5®c]q��!HB��?|��[/�{nrb�J"��ޒY�Y����a�$+ԍqe��"9�G����<)��Xxa�/�(�����8p+���xi��-"&$�����:�<�eI<He�W�}&�P�b��̯�q5?2�r��*rþ �������n�C'Į(L$��e�
ډ������vF���j=Tٶ��	\�S�����P�Кz��O�JW������=����q� �7$Txt�SB.N1�J�z �:<T�&�3�C�ށ	��:-�]����7�5��+��������+�������&3��қ`:F� �PZVy���>�j^j��֠�ڧ	\mg�|�$�������'	�^�� ��z(K���$QI�h��e�@��p?V����vqU�ܒ�-��bS!$ɚ�����n�u%	�E>�CG'�M� =�iS@�E�u�M���5Zј��t�/��*��0W�� ����eQ�?�"~.h��jm(}L\�M�(�5��u���4K���.����V�&.�Q�Q]��6Qz^�K7/�v� Z}�w��M��1�6o��b�8��j��|�8���G��m��r��,ծX����]��CY�|�k� �^�k{�9	�k�sZ�_"DOJ���1�ujYS"z�b�E����a�j��������O��o������m�E����墠�B��Ĺ��V�gۜ^b�;����n?k:�\??�g��+3^��Xwc:�s�R�!��з�od����W�j�P��Q/fe�er�����#�+^D�d-�yTL��h��3z54�Ӱ�x�@?cw�X���t��f؉(�U��Ox��O��`2�K��,a�i*��]������}��%[�^����}ǣnH�_!�t�8�J^}m*��*H�wq/Qf���<�nma~Ɠ\��ǵ��7�#��"��긗��DWݿ���`܁p��Q6��PZ%�M�&X;����A�wl���a���䐈''Krr��6e�)�/�pY�*�D̏�\�uiE�/�Q��D
�90��l�=�v�#Z�Ͷ(Ŷ2���Dh�Ћ-n/F,J%�o;��>��*��r�߬�Gڲ���DO=#�e��%��o릗��Z}���eq�����c�@��&e�2�Ԯ��IX"Î}��ghK[�aE'0��{`�l�(��x���P�~N+$��B���	ѵ���E���]	�J���M�+��s��#�@�gi��<!��E^�<�\�8+�,e�-����P�m�z��[&�/�&���S��1jŏ�f��!��b����xc�,�Yg�V���o�CXB3|�5����t!�~G���o�x"3��\�n1��M�M���Z�}����M�?��)�������M%"�M�{Y��Ew�Gr��@rn{�3d�:���m�_���G��l�O.���� ���7�)��8R��y.wRq��`�W���rk���-7f$l�O��+y�K��X��΍+;k�r�%�	�F��e�e��Sy"�z9A�_��1��ayN컩�,6���	F
��.��cuD��ȴ�Jk�(�^<�$�l&Ml���>!����$�s�|�Ur
���R��VG�z��Jh0�[�J�k�wMm4z�l7T�b���(��E0+ˢ��bͤ�3��k�j�7��?�b���b�K�FPҝC�ή�]��]!t�s����%��	�Z���&h�E��g���u���{�<#��B$�}�XB�__ݱ4Nu�<ŧ̬��U�1���ޥ�q�n�ȳ�s�}�G�ɰp�b`��P%|S�{i��w*VI�t�t�����S��69�ģ�����n��7�E<>#׾pZ��� �m&lF���eO�D�D�O߳S�e%N�{�Y��P�%*U ,�������s� ��w��
����e簥"��:�Q���c5�6M[�C���SeL�q���~EX��nȍK�pnu#U��dO�����k�<+.Wަ�_�C=��s^\�9r�/JF2���33@ݯJxyf�hq���{��.k�r�(Ԃ�¬Ap�`�`�2�!@�퍧O;�w�hiM%��2���1pg��q	[�"��8�ЫZ�GKƑ%��m�~�4#��>�~��g�m>@}AW�o�KT�C	����ǠNԑ� �&��М]���^%����	����k�Q^]5� �b��B�@�2��P�g�V�a����Y����u�!��W�A}���GA��v��m7��I*���N-g�9f_�y�3���P.�]ėm"M]G6�!gZ~ZRU�"�Y���N͔���o'�/���>����F�O}�'5������JNQ��r*��/��nP�,sXD�t�MضkNܢGq7iTyH���3le�kQR���d�;��^�8%�Y#�׊���f���Lk��W��[l-���L]>6u|���B�x �K~���E)�'�J�0�Sg�g^&ȁH�MӬ���C^���P�:�9`�A���du�&���¡���*Z�l�#�J�3����]X��K�Q�� fVM��D.���0 5x~�6�<���D���E�����-��F����몿�ue������P|E۶�����+��5Q��F�&O�^��ribe������,�О+�(���t!5��,��'\cZ��RL��z�v�~�, h�����	�u�>�_;�J $Ms5��i2_Տ�O+���������ⱖ��B<��}%���������������zJM������J�N��������!�b�x�,���Xë9����/�H��̓
�$N!�/z�k��.�T^x�/��
|����]YC�	�~���ib�z�Cת�eV�4^��L�oRͧ�2tC�È�$�ݟ�w@]��
v��۠X9t"F�Z]�L:$�n!�o(�������"-J��� ��E����U�wn>$�m]v���
�k�	X@��F��!�<PJ� �jk�V�pB*i6T,��c�b��o�l��c�V��xN1Pg�o"d�T�	��]Ӄ=~̞ V��C՞�]���-r9������zr'~��mG��m�F�>F�%�*�m��u"��1��QQ$����Û�T`#Y����[�q��D�X�Vg�4m��
%�@�s�kY���]�����J�x=�j���j-�W?�u�ĸ�Dgߛ�N�w!/��p��TS��=hqo�Ӣ�lq���p?��@��)�#���cW
ᦑ4��%�{�Wf�sS���7���HN���J,1�xHZ(=	$ �߲#����LM"Ekk۰��H�޼�>���z���t���ѲB�V����E.)d�
��o�E2�t�r�[�`HD����
,9�����������G����z�x6npƁc����ʄ��i"^�v��i��y$��9�S(��9"��ܩX�i���*��1��)g^�8c���*�g&��iN c�f�@?�!݃����X��)3��T�������pV'����﮾/�\�C����$��D����h.8�G{���Z���믷�,b$��b�]y��F4+�����)?�Gf�<�����[����RL���A�Y��F�?9���Q��\�!*�U��|�O�G��s
|=s�m,4V&����Wv����(_+�E�ޒ~���}c��Dikզ�(Ѣj���� �ןaظ.R��P&�<����R��n!Kd�\K��rL�^�p�l#�-�F�h����tk����s1�|h�T��"�(�zO�Jm��
ș�eYw�~e�����z<Y��;�{��+|jH��0�n�|4��&w�=����^'�i5����ա��R%��W }I���\"� _�w�&�nZ��_,
12�kQ���m���4d�"����������~v�z�woʯSq�?���Y�Y+$2o�(U�%�6�p���,u�H������ቊz�_.�i�4��M��g��7?��L��q��̒�'��jn4,1���$�So��ˁRr�����S^�v�!����y��2�G�S	�G�,������<7Lb8���I�\xU�q��f��1��	�l�e,�cOפZW2.9�G'F�$#��8���(������\zr��6�r����{K��kV��̊� ��7���+��!�q��tD�p�='1Zr���]֘��P�����~O�t��X$��+n�E���l�F�d^����ZФ��Ȓ@�"
u�
e���k"�@��B��J��6�pfr]fP<T1�Gi��~������-���#�K�	ft)ٱ�v �,��>ݖ���T ��!�ն�VSd6�Hb�=W�D�������-8֔���"��ق�i�*��,T�������%�Z.n^ߥu�cS)�\Re���٪��m�Ӆ���x)W㇠H���vNُ��q?�S�f�
�CA��1o5��Lu���i|�]x�ފs-^.�z ��i�@z�d�G��-���+xa6'�ޥ�.���/a~`i̳��(�L$�-y't��k�iq�f<N�Iꬼn���W��ɹw����(�TV����`l��D�#���)wQ�l7������tH�w޵�f�S�Bra;��"a8,Z�nqt:��7x�=�$"�7�W-�iL�GzTmTquQ��]���`>��N��p;	��IT��Y�4�_���T�I����x8����
?=��#mK��ri�3��vUa�)(t�c[XG��V|Ňo�� I�dq���vSo�U'm�(^��c:YQ���Yc���n��$�(��!��AOzَ��0���]Kt��h�.ű��ʻ�������L�_�M[9��.��+K-%��1���3#`�ȶIbۚ��7��d��^��Y�DNnU���+G���y��󽃂z�a����2Z�a�Yt�-[Wy7�}���m�$d����W�3��f��|�k ���r	��[�}T�iR&ɲ@�i���ɠ�>�o�r=�ZX�;�f��??���"���m7{���ؑS�^T�P�: �o�WR!X�W}MqVtʇg�{Z�%]e�@5�]������ �^~���Z��EOM
�-	��g?M��h��z���G�'��4��?�!�D:��$c~�
�(�cI�%�>6'� �ژ�4�$�M�������B|�\ Ht��#�8�6���B'i�^��j�S���CQ��淞���s/�YL\����@]Q�	<5=S@�`�;h��v��Jt�u'�8�b�Y�'�?8�u��U�=��DC�5x��`��.���:��핏8�YXa���LV*���mp�������Zؼ����;k+x-^�����y'`���s�.��U}�����~h�{w$��&#���6ak-I3($^4�6'��:�����"�]����{>}���-:��(v�aY�Ms�Q����Ъ�Va[Bu��~��#���I�k�,���;����B�ة��T>�mmᑷ8C q�@*�AN������\_?j*�^�򥻏�d3̸�Н��ֱ6
߭�s��'w		��۸��kҙ׹�	J��(v}ؑ�2y  �N�X��l��V��1t�����R�-_�G���Ƕ�k&qW�Tj	���^+����"�Z#��ǯ��]��	�֫�u��9�E��:B��S�iR������H	��ŭ��82ϩv�:ٙ��F�nE�u$�-�<��SR(��_�r�G;֙-J��9[�4u���vB/��Խ[��}�� u��-(���XUh�c��I���#dg�G��L�Lz2�wJ���'�^�>YGQc����Q�'�W�Y㞊�X{�=V-�W�8�b�Q�,���ɶ�-��-��ǙZ�_�+sk�G�������5b���Z8v��������G������9�0���dS�{}if�d�k� �P)�'�Qf|����+�,ǐ����~��B�N��3�ʆz�
K{T�m�QXsa�U\��/���92+ q�O��5�. ��A:zf����r�(�Yy4|��%d���"�M㉋�5�����$od��=O��am?�V^=Qr>` t ͌��\k���+C�>8�� =c�������a`j����`\>��$�R�����lnSK�6���J��
�5Lvj�]�s�j^
��p�[��ǳ<H�e���K���o�Y���N�w��j�q!xa�NS�͙<�����QT܋jQHڼ��/���C�{3)`�Q@!��!�K�L��9�
P:>u:T������:����Xp�ų��{~�F*+�1+�k�;�C�$�q�5�ӳ�U�VC�#Mo!p>��Z?#6~6�;��Oi0�)h1t�sk���[�<�G6d���,��A�p]��J�[h@��^�c��o;|3��	_�AAAi��<�@�h��>0�COq��V`�H�v�,~�;�]���Bg=|��J�.$0�yQMtSSmj\�w���^�s��ק��x�#�T<;�
���:��%�ށ���)|���$�.	��n����/hA�[������b��㨬n��Eb�c����Lj�k;[��]iQ�S%TԦ=		�d9���c`���
�4Rt)�~t�Eh������W!�p��z:�s��J��,$�/�.�z-�T�Ӵ���?�,,^��� L�l�jeL�	������?E��	ȟnuI@[2��0X��3�f5��{AC�����fRX,.��T�L����gi3%���+���V��oC��(cy�/��8�u{��ҡ|p�.���O��'|���E��K�È�jFA�����2��K|��e�H�{�P�J�vC4�I��TļY��O�P]qz���w����Ѩ��>#���<f�g:\/�J8`m o�}���
y��SdMD�ߞ<�)
�B<D���a0�)OLת�9�܏I��ƱA�k8{�h]'v7��m3h��U���	R�%K�پBR A{��7��.��=�#�#��N!��Y�-�|f�Q�i�5A�Y�gp�B��ʺ��v��+:?Y˽뙞m���ʂ%��L�M;�;��@Z' �3@V�� ܕ�஢�A�m 1�,-b��'���S�ЂX��]�.����߼ �5��ViFa�$��>���ǯ��-$SA�4���I_��`�$���`D	vc��r�^�,K���O{f��O�zD9h��<�(����4�qFj	�w#�b�4xlt��Ƞz`���=&/0�t A�2߻F�	A�yUh%m��Ù�A���,���mJg%�S`�)�N�]��6+(���,��܏���6A\�%��͞A;��Ag�\�r�H�`�pY�Md�؊-��o��K�۳�h+��6�'���:N��w9%���W2"Qo�Q�,@Uu�2D`㋴̕��ȜRޖ���.ʠ̇�`�������d�ŽKd�#�Ԋ��(R�WJ%*�����d����j!��zwZ!i�w���م8�y���4"tB
�J-D�@^!	c^3���������<Z.����C�;��Vǜ�%}E���;c,�H�a�l2�#4��I՚�� Q��ηO���8�Б_�zZ�q�o<?�oP-n����p!������?q|ds�pB���*�A��s��(�y16��9���Cgkt�s��KV�����������͔��\�@t�T������&� �S9�߲���^��<�C9mH���Ot�Žj�n4�!�z`���*'h���ֽ2N�� ��%�lU�VB?<�[Q LK�$R���/�hh%ɹ�bcyR�g��ı���$!F�.a؈���
n�/Y����k��wν���0�HC5�?���l��ǨR}��Q_8�jN�std�B�%]��n����#��&�bq�������S�V��k��ޒ,iDI��nq�yP ����[���oR���Ձ����l�گO�e$w����H&����^��8��xSg��g�-j�Q����矬�Y�iL�އ�K�*H{���(ߎ�f���:\%7
���r�!�t�5�P��[��sx�%��T��-�}�������WL�
�������)�%�h��ď��D���1����tlP�ٻc˫��^+|��/��ս�3+�O�j�>xk�.�t�֕;ĸ4k�k��ݯP\jkG�S���Y/�J^��<η	�<�+=��˘�b{�b���D�h�{�t��۪�y�6iC2�`T�1���^N�FGvh+:��R�n��n��l;����2;�c5B��	�oη\*��w�Ϙ�yy푍��:�^�\�^�V�%��Y����� 6�U��u�s�P	��zBM�Wq�o�X��bZL��Y}?��5n��R�F���Ì��i�4kk�v����/ֿ�kV�}�lB�� W�K����t�a���ͮ��-���s_���9��b/�|����it�	��J����x���J��������߱�i�*B���L���x�	�5 %D�3n��t
7����� �����D9*V=�|�s��1i7x�������n�)#��4&i^5�n�R�r+��{7��-�RMz3�c*A v2n?{nU�L���'t�i��	"'�M��X� �Y��Y��������[�`E	���Q1z�n:�Gb�[��E��� ���g_��{�R� Z��f}+%M�f+8{|�sB�����]�k�[�	��4��\����ڎ�����Vؓ@?�>e�CDI7�	I�R����A�a:���!MD�(�SD��K��G)���HP�S�g�GLeB7�4*���}�7t�������~K7���!�'
�O$j�&�a��Km������SY��=�M���#�ЗDwZ0K��@����㖵J¥�W����25{1u�!-�1 2�B�_��*�]4K)���3����Y֚p��W�}�@9U륥pY�.s;N�p�Ð��@_u�̪� ��	Fi�,j̢3��Z�6�����4�λIF3~E��9լ\�p�#�${��ʿ�ҤT<l��S	���%���[yB�d����}�hS��o�>k������aύ>(� ��8����Y_@K�e�pܼ�e����9�b�TLz(�ۖy&�#�9��w�t�eH�9�!�`YWQ����ˍ�a�dQ��1(�.e�����\w`�WU�s�⁠
J�i�í�I�;40��Թ��ek�p"t�V���>�(�E"�`ň`�S�[��1�uӻ1'�J @~��z���ɡ��͟�nk�W��/�|�^����]f8ߠ��o9z9W��F���܍��H�
^x��5�Z!�@N��ۇ�@/�%֤78�V�|F�y\�@zW��w)������ǔ��1��A�^%���Jl�h�s`W�	�l&G��7�0��΁�v�̇Uik�9���Ǘ3j�{��F"\�@��5�p;�����M�l�r]����*�Δ��������ﻢlU\��=L(U�3�\
6��1cyBYp��̓�ǀc&�<��`��o}�!����k��۲.A�'4{oc�P�=M*�/� [��#=���{tz�M=<����X�8	��qE��y�UFD��0jp+��5H	)�'��"�KJc�p��@��o�,�w�п�oT��&����!�������xB5�rQ�w<0��b�_��w[� l&��7�C\کdZ�a_���Y��w�9w��.�i9�ӡh*��l���W|C���f.MfR����2�_���$w���d��}C������&5�|HK|�M@/"�L�F��G	�QE�*9aI	��j;?�#KE����EW����G������~�,W�X�����\~�짜W����⠬As�o8Ng�%E2ʾ�@8zEk����w_��`�c�{�%Oo��ڏ�І�0�:��[,��=��gbUJ@��Ħ��C��0����8�7Њ۝J&c� k՞�+�h�*�����@����y5�i�~�>cc7ⶊ����S]�V�����������x�.�ޟ+�uxN��S��B��v/k��hM���v4�*�ڴ�|^lSO��{<�"�x��t�	�ʥ����n��j')��T$��1�2�>p*~q5�g��� Ϯ��^�C�����s�KX�������8�b\,�m�_�łJJ\�ߎX�Z�R���nB�+�+ma���
�E@�c9�se�:ɬ�`ٷ�K�74:̬��n��h�xc�/�R� xĳ�Q`�6�K�T�(�,��5+�@J�8� -��?�H�fR@Br5��4�2��h�䥣m-1m�L�A��y�4i���\��y�X�b�׳�yx��V��/���o�j� �8+B�r'3��'.��,yƉ ���n�
��X#ڄAf�:��]!6$���q���߻/{��2���RN�#1jbe��H# ��Tc�YQ�O�M�w�9��Ŕ���\�>ө3eM� 0vțJ,����o܅?���!�[ybD*}㓛��?m���۽�ܪ���4ů���+B��z�I�}Z�	t��zu#�9���s��kq�$[�� Xs���՜�3��4o}�܌��õ�����M(�U%�kן�����vVZ�e�u�1���8��[$�2I���
��$��2�.���ME��v�}5x�p���>�Z���i�*�Q5��h�4�/j��<����m�&� l��'�H.=��"���e�+fp�ၫOz�c���2�n���@���y�推�3����LY`e��aح��Z�����'�Mu&�1�l�XLrd���2�d����~J��d�*^[��=�w�u��4�/$t��d$�(S,ȿi��;m�!�r��rX_q�g-��`	��2q�m����c����)8Y���3Y%nl�)U6� �9�Л¨��U
ǻ�A�z���~��}A�B�
�т�n%c`]3�,>�%�I�C�x�*���|�pm�n]Ky�sn���_Q�.^ţ�M`�Q�ց��XW^K��iE]��U�6�k;p���R�KJo�~��5ڭj VH��j
� j�F��9�%��?��o{��Ĝ���*��
�w�ȴy��-f%�t,{/��Ȇ�܈���,�t���j@��г��lW��FH�M%���f�2��=Y
�J�◲t���	:���n�-;�d}��U����Sl6���3TO(2l�-[���Ћ({�p���q!$Ҧy���A��ġ[.�����Y����Q�.�SXT�S[��3�J5�}8ߤ�Zkܷ����u9�7�E>�����B�X]��Q��%���8�]J8��r���R\��Q-*��Pޫ� a&I�<�L;o�ˆ��c�k5�}b,���=���^��mT�G�:_g��Do��E���h $��m(96U7��wV�^
C��u0���*�n�"�tT3�A݈�P��n�� ��s�iK�a�fP����
�P#5Zp�b�y���.=w�1���$���\HV�W:���� ���q�Q���5��V�R�y@����<�I�e>�����֔1j�T���!K���ն����Ү������� ����y�IO��W?ut�gP?ba HЮTC�֩��'�z�Ŗ�O�33�����=U���i�c�D�B�N9d}�*���c?�^����7ߩ�S*�AViɦ�����zW'������ߓd�-��܌���ng�Y��%���S��B����K�T��lke?�5'��m�Q�����
�A��?��Lm����V&i��>"㯚�s�.���R�&l��٭��ec~�ͥp!�u��*}Δu;g����#����5[%9�d��g������E�nI����k{��X_�`?�$��:����p� �1c�$JqZ����p�����=	�D�A��kFH"w�S�w?7ɻ��V��՗8r��� ��[�jZY����	�Bul,�(�sn,�'Vk3�c��<HC��w䴜2lq\>�ټG��\��M $s�0����ҎA��Up;��x�t�I��h�����M=�o�2YZF�R�,p������0��SzG�G��Z��x��ߩ��K�4��G��g\��
��܄� ��@�Nd� 1����?�4���k���;�pq�D���8���Zp�,�I�2��j�&�|M;V�ہC����W��8���\�hc�� �+���5��ǎ��/�e���b�yM�)�J �X6�
�U���X�Gy��R���D�u������Y�`�3�q��ev�l��������.)�^�<�?�P��M����uah�:�#�	��ɩH��H��0��?-��^��	�[�6�����햟�[�5�F��r<�ɡ;�vq��q�1�=-�u���.���&���!M
�!�G�^�fUr�:�Z90�� �Oܮ��1_��{@��sx�_�=���r�L���lH0��Q�&���A����,�(���݀� �#Y&x�hL�U3d�i�$��B�r;\���1�Yw�f�dJ��g�̞���
O�Q�.?beX�g@-�ƺb o*RGB���q��2�)]>��.&��dL{����u<jn��	��du}�V������)����6&,)(m�o;��6��������zI��A��Tz4���3�$����me����Qt)*�(9_ђ�Y/�&9�gWa[o�> -]fSJZ�:�_4�VE��e_�r��ďm*N$+�[�]Q�u�Xf�;�UO��G/Ҿ�b�v&P��;f�1%+��U���a54��3g/�0��|��Uw�o��P����&�t�>�.�-��������*�n�/��+f���	KU3�'�ס���8&�z$���[B���`�Ww���ݰ}���(������WҊd98%� ����c�g��t����uBP�q�,�2�cYN#�����[�8M�?��[QH۠:����LuO�$���6��T����G[��v#iE8 �7N�����mQꕕ�H�}�y�8���ܔ/��	n.�/�T@iG�,Nw������J�j�6�?���%�n��Wi��1�6w�wJ(g���ECyG�CJ��c�������ZH��pTo����W����	�`����1�A���rE��C-�Q��q�m}I6I�o���$��%��e]H�>�����*���jJ�����Bjz�ڱ�6)_�_���69Q���K���vgp�;�f�W�s�{=��7��,|���Iq2�Q4g��\�uK�hF�h�T�$��ޓ3YO�`;���s�pknG8��˯�[�"���.zV��la�
�O� 'ᜡ2��7���� /��\�f��r�$�L�"�2�n���N�a�I��k*<k\i$>˦�Q�R`s_�H�#��A�so�^�9ֆ�+�������.syvl��u�M��H��U�liD��W�l�WR�4����t���򆚛G6${ZƅA��X·YRJ.��l)Ð�Y����l
�1V��k�OF嬬$B���7S!�iU�Y��h�p`86�-�ԏ��Q3���r��A��#R�A�����W�d�XmA'g���(���w��й�h �g�?דE���[y�..��X�����m����Xo�����҃!�.1�y�8{�s|ۅxtóɨcͽ��P�LV\��^��!��s$�,5+�֑N�&ȵ���h�]�)�2�T[��%�^�ۤ�w<�� 'tz��B2G��:���Rs �����c�"x������J	<㇯��kh��h��`)��H�+�-�!Pw �����ʙE7��})�$GN�GCQ(��Nyэ�=�ѡu��2���ծ��ydGҞ�Z�ZU�m��kFE/!g��Sbf�`4i	�-Aһ�­k:ݫ�I��/��h@K��S��*\HUQ���Z5���uDJ��7��ߊ�"���h��L{�#��W�ܑ�@>�;	}iw~�?^�_y� )1~����%[Z���Ě�o[�����<���<�7JՎ�_�o<����)7�݁��6�J��EF�y��.�z�6搔Y�KƘ7livP��N��ʘ%��s�
��0Ǩ3�]gTK��bH�~^�xQz���O�T60O�Yya����h�6_��Ӈ;nbY�����JJ@��c���-�C>d�%���L]����/$��9|���u.���:;��D(�6$�����y�$�"�����/��ڏ�I�H�a��C�SL(%�_ ��Gμ$%39x���^@�~!Y"�f�#r<v#�4}!�<lܹݲ�����Lb!�[��h1+��c�)1�&�G�yT��\���.Ga�Nr�}��H���R딎��F�l"��Ǒ��>�����]x�X�k̊S15`bwm����J)�T]�X�31*���PR��#�"�ȱ�ž.�3���{[�XGr��`��"QkG2K�.��L)�P��3�4���>�0�{�$��Z�!������Z��%?�����U��Χ��[�0���)��#r�q$2Bl�'�I_/����ےߘ�|�q���N�}J���D_#�/4���P���1ZY��
 �	{c��G^ڵ���4A!و/�)� �����i*������2��0�_�֟�[4Սѥ���HB���Rue�˰�%�6��p�����7u<WFSW�T���;�l(�N����� �{�����h�=p� ���ஷ�����@��:պ�����}�D<�7��D^%�'(��ӏ���=�����_�Yer?6��"t�j~g;1��.n�F�9�Œ�<����hk�p?�^���$�.ឥ۞��[<�,<�hj@)�q����_|��r%���C��DvB+	uQ�g�ѫ5Z��ǵY�=��Z�_�M��^��(�]b�Y�،!���Ѻ|�M��.��)|���̳�T�H���۬b���CGE<|��7r�{i4�E����"�%��puӭi��C;+�ޱ�-���@�怞����Q�3Z��1�\d t=+�ѱ��W���\�keҡ�eUaEk�>��MYf��������m-�� �9��)�9�2�t�+^�i����M�)��N<\u��rE�7~
��Sh�DL�0u�Z��'\ �0om���8I���۾�n�y�̕�;��v�����ˊ�m8����4� ٺ���b||� @[K�mxZ;�L��)8A�
�ڮ+�m�x^^f͢L�ǘ(6ڈN��Tq�Y���lR}�|*Aa�{��avgة�dB��w���<&Cc	?���W�.�]�}j��4'�k��O&���ƛ�m��\�4 D�3�)?�|�	}mK���Hsۖ>/l�����;����'+�@����0��\�D����Ti%��G��u �]�1���D�n��p��w���U���=!`�������ځ���^.֩�xYLIL�o�"Kf�ԍ4�����K�bE�f&�D��{zۢ�I��(��v��c�r��j<�k�����a|uY���^`�V͡;G{��8���W�2G����0e�&Ti�l����Qp��W��u~�tK�C�����n���T
)�Z얇4>O�Ķ�'����{�z}U��V����a�,L�V�)�]o�Δ�o�����s�.�Ut޹!��YL3��6$F2�)>�$�J�]����G��YnFDG%�/����J�Q�B22<�6k�q��k�����|��3N�w�Or�}�2��?��벸I�%�e�Vk3�bgݷ�(^V�Y/��p���9{L��^���дq�m�.[�<��}jF�v����zY-g�'֔�Z�o!���#
8�0�[��@P�~Z��g�L�_����*��V�e
Mɲ�gVk����F��<J$�?���x�ڈ�!��_p�b����v�jN�	��!I��,!7�<A�%�!9�j��Ff_�J����V��aNZ/���}� )�՜�#�w�>y����<�Ǜ��=�頉~����i��b4"�q������u�i �BMOOBð�j;�J����΄N�VHvD� DC�J��|$�C���3(ҽ�/�<Y_/[QBs�K��|�ꍬ���羪�Tb�_��γ��I��IEr��geln�D�}�4�uI�Ұ��~���f̛������ ��X^�Sd��7��(�d�Sm�P#ℝ���L1k���̸���7R��4� k��� g��+��t�U��#sf�0������u��ZH�q@�ra�t��&��A!ϴ��גsB�'�Ncj7�Z��ʬ8�kM�:Bێ�!��W˧;ngf��]�'�R��.�]�k�;"�6��t�����9\5��
e�uM�X]
��6#�c�ꨐ�>�{8Հ���Lu���m(�V��qY�^���ܔ�5Ev��a�ꗞE�x��j�P�8P%�q�v�����f����-�į�7mZ�gT�Q21إӔS�o"�pv�M$�]��-h/y�y˹#���)p!��?�Ē����"3�+Ѷ��7���.)웫��T;,���w�D���RJ
S�j�W+�_g����.�pC��ƣ�TUSs2�O���|�������j��ݫ6�L�
K�K�����hK��"P�=1������MYA0��:�H��\�W��� �Zzn�YD�&��<~A�����< #��8vkJ�:6����y(Nk�m�q�C�5K����r�}{�E�� u0���>n�jX�~��R������z�A 3�x|A.�t��|�	�¸��79��}+}��T�z��@�6�34P�@U#�j�-5��h�205q�_ZZ�0{T�	��[|��y� )u2�q5�H'�|���|�����͕��,����Mc��
���<���5
FfA�����o��Q > wd>����_NԺ�0
���<�䉻�u",���@�i�K&��'�Iɽ��vr^�ϖ ���1����&���ܑȭ��7MnCĠ�iN���Sp��~̓oAlE���\��+t�z�˓����z�}+g9����㫇1�ݵU��#v�9�3e����&�Y53Y�pA�� ���U��{�"�xr)\+k�{���R��"V4��e��CH��Ӡ7�S*E3�SK_�E�_�1��3?E�N�&��ə����1Ip�H_mw�	��d wƞ+5=��틊�{T��]0�`ܰ,tB]��P�k�q��f�i_�Q-�����a�h�a�;��m!z���4}�
d���	D�(��<��y���q�a���zCU�����\ؒ�Q?	If������Qw˭�<|5�g�'# �7��Z�δ��f:��w��fo��\k�lGH������T��0�0o��_���V� ��Cj_>�TrC��k�����/�D׬G|�5)(,�;����/�ɐV��]�x˗����}!J�K��� ��xdj�%�3��"�y�� <��
���9H�
��{ÈG�8n֞|y�=_�^5�Me{�X�C�@�e��c��CWNA�5#�7+G���͙d�15���W��c ���C�*��A9��o+�J�wt��%�{��j�"�"	�8�[����*�NF�	�����@H	�|I�����ZƵڊu��A���d�i�_��['Z��C<�I+'�䀼�U>�T���!��C�{EyE��xV^-e�?�0�N���3U�y�D+s����˔AdnT��ש*UN���^���}ё��X-!�1#�L�1,Qf7u��|W0�!�rT����kQ�@�,9�p�X8Wݨz<��}�@m�5 x��uld��j0��|<K࿤�����D�8��d�kuȡz�_����D��̊� �(�I3�3~��!l�_Lw��T��c�g�">�m�"v_ ����?���Y�����NC���,"������.¤��Ix�q�!��7Dcz^�����<#�dx���6�,�x�y!��J��t$i�٠�� �Zn������}=r����1�%P�KFU�R��Tl�h��2�.I@م�� I�)��n�zB�m��E��G�jJn��u������Ds���2}6Do�܀���)OE.}���ӌb��Eİw V���G���J$�1���z��[��sK�aT�Zi9sŌw�>�8p2B�I���K������X��ƕ��fS�^����h�#]f���^"��2k��Ox�9\�~��C���#����=N����m�4����G!_ެTN��~m�G�\vu��k�u��W͓�;�n�=�[�>�6	Iϑ=/�Q=��s��G�������Uf��&���Q���,�!��W����Ci�$�%���9��'�;������V��0d�g�0:"͵���UR	Q�u{ӊ�5�2d�0k��X���
���P������e�O۹�7����Ӧx&qɹ�j�5hN�`�Zdk�!���܋|�5+�����U���i�����4��`E*�~�;�v����e{dhWϘ
�ϥ���z�B rw� �����n>o1Qk�4t.�h�T��8�����6�Q�'��:l(d@��D
.^�=��kĉb/'�ԇO��Y��`rQǡ��7&�	�C���h�#��ʦ�aG�r|�����j��m�Q� ��z��(�Q����cTQ�j����P&6h���XxFH�u\o	t�n��E��^6!y�*��0ۑH�b���,�|;]�6�d�-��t���a����>`3��`��Txђ����{!�m ��=�0w;"����ۈ�&���\���ՙ���W�VA�Q"ͨAI�<P:�׳���������w�O,4���G\�e�e�
Y��ь�<��&�`�'�Ґ�.�(�%��k�wh�wMW%UTj�6��AW42�@�jp�B�h����'�^Bo�Z����K�'���?	t2�
��$��1*�ͰHi#p�7���������|"?�'�\���61e�r��8�"(5�m���$�5]�Nz)��锩����6���"(1�-�ڥZqte5��n7���4sAXr�H��i��KL%�&�k��f�]���s�3�ZYo�!s����~�x�X{�PjY;?�߄G���8�{Z�ꋷ������su��	SO]S�z������0�U�}d��Y���Dj|㚄�њ�����(�Ȭkq��ʻ`�#���ɹ ��xyȃF��[X�׿քb BN�r�S(��D�s��<��`��ҏy%������N�_N���UƮU��烊�Dh�8Y�n���[j�k��Ǩ.��Ź<~���= �F�7��U �學����+uWPl-
��$�K�[��pJD*jp9\3.�z"PI�vW_ۭFi��G�۱wː?s��C��}2�J��X+y|�z��9x-�2���)l�=��"�
�:�;E�(,�@K�\l�d���D*��3Ֆ-z�>����\���4׌aT}��X��A����'j���pO��F�e#b1JD����!pU�#"��Uk.�(�!i�TqN���{����C�u���^���р���b�v�yp�Y@:&:Ww�2Є_e����Q���B*��L���>�߷��a�u�o�?#��;������r��r�vYD�FD1���j����b�s�*����A�~	��(uf�{13��D�R���ڽ�M��Qx���#5 &�獒ɩ�봂��~��\K����"m����|����
Y�CHu�����F.�ļ3~�b�;�ztCDW�<x�d`�yԈ�^g;��s���R�bj�F��$.�0�{V޲��s�)p�<����hY�"�)����W
a��C�˨ms~���7�[��+����˽�׆[�G�o%�2�鍳K�c�����yuL{�kL��]$�w�C�՟v�V�m�,P<��hO���,3@B�Lb�>Kkc����}��l&�##� 68��/ZX���XE�H�2�G&F�K�F�P0J�`tk]��Z](�6���t��d���]|�1vS=z6u�Z&�R�MX�-��-�КH�o�a�V"Z^���NT�I����kZ>�� �D��[b\BE�龶@j �������>���hd)�~����XĿ;oD"!�|��J˺>�r�P�)���*O;�H�xٚj��ʥF�X9���A�ks�ܜ �z&w7	s%Umq(m�f
i�M)�k�Lf�#�Q��b��!�v���(s7����ء�����N�~̐rln����$I��渡۰����+]�-+�G[`�$�YE�QV�u6g��xB0��<���� n��LW�.�[���������Iᗺ��W��ϓ��a�R/�48V���$i�'5�����V��ކ�豷sz{_���v{~�]׹���ɴW�Vl�`
�|>D5E
t��&��h�z�Èmb�^>�N=�n�����)&��V�n��[�*�*s�r��.u̫�U��Ѩx�j�3w|*���F߮����ͅ'��~w���X��F��,<VL�>�lD�K�M�t&�\fW*Iv��tm?F�s�	�N��0n�H.��<�X�M�gs�߮(i������nH�h���)�O�;��K����(�HyyO���j�Yx�ݘH�M̜����7ɣ~��v; @����DM^��}��2�f���E�aĩ��V�姦�Xԟ�ӓ���Wكt���\���"��b��+��[�(Z�:U�/��J��ى���䂀>�B�7T��G-�����loU(i�SJ�4��*z��aީ��Aȳ9�lg��H���ڱ�OAW��!\��^�8�WC���T,���JH���/���n��%��[I��l��i���L�}|�R�R\��Ƌ ��1�2�Y�*j���t�l$�-]ĥZ��K���\�;V۾,�F������nۭ��WN� �$G�|)`U/�����P��4�!�r�Qw���S7�k嘔r��@*�T�Ɵ]�Io�/�[������������ϝ�������#��D������*�˗鶋6h*���na�<?�x��Ho�;�ZOTJ'U��G�nH2��k2��$^+�f��~�H ��y��4K@f�h}�Q@{�!�aj�JV#4��x5���TIJ��=+'l'Vbx߾_�pE��;>V��.�7�Y���FB�4
N���������.C�M�Y�aC����t���!jtF�7����\ �;˭ ��ӄ�W`�ڐ��T�)"�3j1��R<�R,�T�_�Aq�M� B����X�\�CtAS�5�F�,|ɳ�W��4LK���z-O��k9M�J<Y��EڙU�^)��g�g]�v�ˌ��[��׳�#o3��2#��f�s&��0� �"�gS0�7I�����q~$o������С����b�;T��]OV�ŝ�y����(p�Gǥv���D�G*e�ЏGvӡ �D�Ҳiqf��խ�xo_w��Y��}�a���;��������O��U$N���_j�}�g`����w�^��x��CT"����D��ݕc�ʊ��`H�|�+O�����T�����YO
�ˋ��[��z�Pz^��挈p�N��h�t�'�,�\�%�H��t�O0��@������\�6�Ƽ_�,H�X��^f2P� �"����#��;�÷ ɖhㇼ0�Ky��]E�Qd9�w��r��j��r��h���%M)�A� ���pK�Ἔ��+���k $��*��E�o�q�q�����ɕ$��ݧ��+%ک������s���td3�h#����C�0̗�lA�i�ۏͨ`�.PQ�)t��Y���'�Nڷ<Z:HS���@�rE�v�G ���e�'���o?��K�����<3'~�7ڇ�dt?�-If`�(����!I� KFP?~a���rA^g��봍WT�_E�3�Mc��@�n>>!�sQ���zr��谔��xv�F 1D	@^�:��"�I��
�p
�'<�Bd��pJ����$�?��.4/.36��O��ue�mǒ2�9݃�e�y@��#w(�c�y: i��zK9���4�!�ET�eH�`��w����>'�/#�W��x�AsvDJ^�=v9��F���W�oìs��2kh�d�B8����������8�t�ʺ�M��"s�X��5�ŢHo�A;�-�Th_CK����I{y��.MՈ� �Y'� ܿue�`��+!<�{_8DL���M���%ݎM�-�.�wќ'���8e�:�e{��Y��m�������m��R�$h��?������pf�n���+Ի��B�X���ńU������׶X�I����f1o�/g�MsW p�$]�4F�F+�px �"j�M BC���{���/���l:Pn��^%���nD���B�}\��j����iK�ux��r_���k�����P�?x[�S�f���X����`�!	Y�H��Z]����A�![l򎿞i��5[x3�p�vd�� �Asj�D*�Vj#�
!��Ļ4k�>���,��F�� �`��~^T���	|����9�$�N.ü�y~��ٲ���PQ�d�0����,4����ѝ�yX�k��o����ӻ��f��4�	O�xD&�H��������v��蟉��CZ�/�[��M����w����@J6�_K(=��jr��%�.��ւmf% ��²��6%
�X�S���L��µ�+��z�1������9|�2�5��_�{6�F&"ϧ�Rz�pvX1��%|��(�*bT������`Z!A��r�a�A�Z_��1��	3DN�g<"�=��1g?p�_�@�L2\,��aX�$��Y�.i�@��俔��̢c �[�dV&�@�����8�Y:aF5��ap{��h�ߒ���8�Û�q�O���^ܠ�z�[%��`u���}�A����@���q
�fb�-�����d�,���~d�V_��ޤ���-�B��3�H�
���a4�;��K�k
������-�\�г���L|��us�>�b�HeI�܍Ճ��I��ni	�w	$�<����Y^�l�R+l��%a���5~ �3�p܆���]�	�8Z���h2��J��BDE�=pOފ�����@d���
[*�ϝ���A[+�L�93gEX�pd��wQ���zr���"z�_٠a�ڲS��+���v��ėG#�F��ѥ���QS��#�]hn:1���a�VYHs���mJQ���
&eم?�f#��1w]��:7G
�
(�_5%�v�|5cB�G+ n�JG&u[3㦥"*@��M��q{���E���<, 	8�?a�mG~֍�b��!
�������F����؅�-6\�%	k���K����D�E��#��8�~��t����t4��L!�oD#��K���P����{g�"7������{ƕ�%���	�,+!Y�H���۠D'i��T:ܽ%���.���OV<*�+��Ѡ�u����=��A7�Zr����oz�,��|�odze�z�ꦻ��^ĭ�{�h�;&�a��dש�'!�g+H/'p�٠�9�����G-�E^�W��з:	R;�B�)O�o����+޸Q�tp/x�P\�ii��d����Ī��dk8
��=حks�Z3[��<������GN��Z�'��z���KQǂ\P�����6�ɢeЇO@<
����)��01����B���?����ȧ�Pa�B&�3^Iu5��J�����O���uS��y@�cY���A�'V���$O�6|ޡ�ڹ�,࣡!(���=����r�V��y��$ �U�z��ʛ:qo;_�!2�jt�5(��U�=m�m2�	8�0�4HXf��r�m[{�?��=W�)"౥����?�}X��q!(� z�M��~��"{�j�EF�f�F�L�RQ�ѯ,@h�$Q?���ll[D�> ���=IR�άT�4������`��:�#/3lA��`��Pr�ςY@5"�3&��0�d*k%����,�Ӣ�]5���T�K�+t)�����fc��|΁,I��[�&��.�����ՉUP�C����nH��.f!~?�ە<�gd��z�:Y��ׯ�)_�֛J���ˉ|�f[
�5�c@��V��\�(�7��r���N��f����ِn�V��w�"�Ȩ�6Xm����<n;+�P��uޒ�ۓ1e��B�`# ٭㹧q�N�$kk�}�ݦ��6�%�v�~�F�|�����a)EJ��>d��ܬKd��>Պ��=Tf~c�2��P�p�� `'Ч�.)���v	�|�X2퀭m �t���;��5�[�|��%��-҃; G��Xb�_�I�Gh�H�ݧdę��g�bq��1{R;�pJ����A�����8+�����@�k���t��T;#���ቷ��O{��b8oC_���by�LGk��V�Q�碐��h�e��})%}D}���Z&��l$�@�	F	7"��n��+Q8��~����t������nk;��;V⬌��k��q��6���e�tu��W���b�zje���ܙ�'���in-�u����F�D�݂i�><x��@8n�r(g���Q�q��W5�s?�Sz�
/�$hY�׬:z�Q�'�A}O֕@]n�J�n��^�]TS��O���r:j�|��l���$|�k����$9��X��Y^ ^�o�.��g�����ѷ �����9P�y��љ�}z�ԋc��3)GMK�E�����k�ӯ��}uəA��-� (2^�Y�N��[o�U1`ĸN(]���kv��|-qW9��R���1�kH�힮�=���e�� ��$�q��7-�gX�CT�n�K!�`���ȑ��v�P�C���S�^hcº��&�ġ��x�ɖ�%��/�l�{I*�m#�, �j�p��������b�6B��������P�7��l�o��d|�������Z9S�a�j�}^��r&q 1�]5La^��<�L g_@/�^�Ҽ��/���-Wэj���C�R���齈��o�6��>=�F�����C\���#�+��W+�\N]&���#�\V�������~�I|�^�l�f1|�����گ���n�$zѴ�g?�J\��e������F�p�ၢ�A=�7Z�M ���n��|�礴?,j�ӎ=r]87R�4ړ^�C��-�?{�x�~Ơ�g~��O�)�C��Nn�[���ʽ�/��61��bM�(�,�"C2���6e�^�".�aC*?%~��5���fFq��M�Q/l�;�~�Q-��3Uw��8T��a&W{MK���Ԗx.�!W3�|�\���Q�5ձ� 5ï��}9��6��C.�W=����X��̌8{b���nF�C���: �G�N�?O���Gw�i]������By� ST	����#6��'��]�R���z�<P&�>�j���"��8�qe��y��j`����U���Je�4�嬉��A��Q�7�g��m�}_�Ld� �9RT�?���XH QD.�CӞ��KB3��j���;��O�C���\���c\k�n ��?�p���������0�p���ƣ�#i�T�Q�yU��- ]�u�����	�qQ�7�"���"�[��[�Y	s�6E�<��^��p/����߮��scC��/��ٲo�/�F�`�Z"���Ƨٹ�R�s�#�@�rѹH�׆D��!�̺#ݝ�]�p���:��gn�Z\.Z�E �r�{��w����_b�M���/3#87�����a���;����8���+nV�)�&]n�yRIY�\�4�&o":�7���o������{�K���c>����Χ�����U0���z��E�Z��.-��7����bNhZ�t�g��mxG���gX!��Ԫ@��h��8����7s��DՆ�q�lp8�=���P���gޥ�YE��.� �w*�(/�
DD�}����y�cn���� ���J[f�'��G�#؝o��g������ݘ�K���9���D$�?2��g�=�Qځ���I���TL�Ň­A	�����f�ɻ�m�pI%'�7�w�/,���+��Bspb�F�4�0�9����夘���?
k�u��~�#ЮRo�X#?�y6��x�_А�z܋�/�Y�BH�D��̺��E7P�6�p���u���4�O�'�6@��75��M�9ȃ �g�A�N���ӓN&k�U�u�	:�,i�;�#�����H6��)���u�_*Nk�h߯�}e�n�S����ţ��7��}�aa��S�~���r�3Ps���S�}�*��f�d4�W<�ᾚ��Lt����F����T�o���C�s���$�p�d(�ف��6b�Oi�vc����@��`����X'rO�:DU8H(&ҧ��p�:r�A�"J-f54'�dL�p]J?-Pb�~���$��?�l:+�%"$��&ƝQ7���zTܵ�����݊�����a�|�c]M6Q�p�~e�1��ǫ�ɑ����v&fw ;G��^���2������Ye��iZ�ú��_��I��<Xc��K6�~������C\4�I�P�6dK㎨$�;��G'!���ny�*v�:e� 
�/Ar�Ts�͒��{�xf��$3º��xҊPg��G�n�����g��_�17.�`�������;��  ���S���E���AW@0at�g��m��S�,�	h�&k����'�{��Z��M�)K�+�ؕ��$��wฯY�pf^�0�9So�Df ������)*��qNL�"���U͒J>5�gBs����eL���΁��md���6���k�>�D]%A����w�T�LDؓH���>��:C�ګ��Y,�p�.]a��������fg��$B`�J��d�V�ׂ��w[H�լ��hk cwnTɡ�>�W=�Ձ�R��4��%�<\=�����p��)���䬊fk`�k��|��5_����FE�WCfFe��Ǌ^��L����XӘg2<��>��Fך��;�t�����}�S��Gі�me��aH�UA�i��X��F�����Dz�@�{�q�t���!��х(�!��^J��Ϛ@����o�(�~訄���F.��ȗgFl����J��V��(��T�/�):��4�2�b-���5�0�\�Msı#H���L��;�]1�ӏ�۳l�%X-1�$֗o�<]���jo����0=�WR��*c�9$�?%:z��x�2��?>V���zk׋ů��-mgL����*-�@�aDy�)Å�YQ��0;���:ỏ���ԗ
3�P_$�7�� �AZ\6���9P�O���$I[	?��Y�;D�w=j�q+����Jkz*���g�%PT��z��7���v?$�P��D^-��'Z��[[���O�r��e;��|��'�g�3�v�no$�����AtҖ��~�8�o[����"��܏x?�<��pD��ɕ���0v,j&��J�£Y;-n*CӖaJ�{hS�"�;v%��&d��|��bטN��D��T�9Ϗ�T��_�h�:Rk�������]��Ö'tj�eEse�0I)7Q�<	�	h���y1��bKl�O�%�%ZJ
/�މ	����dX��aX�% �X���Ji��Uh����rҮ���+�>� �?��f��Kf��2����X�_��௳"�w�z��R}���J����X���+���xo{���[�W�l�CG�����
����)�i7��T��k�)���ߺ��{k'����f������V��s&��a���⊳e�eh��I��
��� l���u�Rp.uF�o'�1!y�?��Fn��,������AX��X���,L`d�!8l5��Ǧ3ѽ����^H*b�֮�nƩ*
1
^�Y��:1t��{jr��-���21�e�x���x�n��7���ﺧM�(��Y�7k�=�[ؿ�a��~,j#qaƢ���*���I���>��~�yc�yd����9���C	_� �y�%6�`><�
���P�IH�������f��[E��� �s҄j�Y+LNml�s��<�6d2���R��㽐�-LH&U���7�;D��_ي`���aL���F.6�p��Vn��ǿ�[����,D�]SļO)6	��/k��8��dRS�� #{��O���C���#�N���%�O{S��ziͅ[ڠU�w�e�{��S8<m�A_�:��r{���9R�q�c��O�f����A�\�~�W�����i�Q�l9YE���%�{���&��M��#�Q�����4 ��Zt�N�y��v�/���Ɏ�F���=������]~rYʛ2w�-��!�'IY�A��(G��7L��hSa�'�3O�5Ȣ��ߤ5:��C��2�:�z�ԁ;����H.U����@�Ja�Iu�܍���FX�ԁ}� ���
��Ԑ�k��N���*��Բ���,���XYee�,܆sw�ȄX���t%�r�o\�C�USV7a7��N�ӽɒ��Ѵ[�窄sM�â΄8��;�-%*���F(���<�J��>�b�c��kQ�d:�����M�7��o�Gk�0�Z���Jx�b�$�Y�<��1X��FRʐ�p�p�f��+.����vt�Eϝ�O�U�jD����x!��H�ʟY��%P�x���aE�WF
�A���1t�̩�.��yJr�����9\4�x��u("b�KBh�W�v�C����O���v+\�7���/�G���ə�Y~�B�J��qs�����t�j3�Ҥ�g���MM�>6g.<Q(�u6�?�9���s����:WN	>|A�jBc��Z��=�.B�� -ncR<	4M�i7��˘�eZd����Z\$��|xó��(E�Q[L�����M�_И��M���P<HG������,K뮮.���������������X�:!ɼ1Q��*-��;�5\J��q�����6���}՟�,�x�6����������m���>r��˘�E��w��@��k�u�oP�3E��j�a��@w3��v߭UݔVJ(i�[a��Qߨ�nO�Jh�����z�gW����EAN��T�$H�J�X1H��i�L=k����
��5���,��|����<=M/2�%zR0-3���:Z�?��H�����ŻJ�l�,��'�ۈ%Z�
�9�k0a�V%�:�h3��k�0����k./Xތ�!qj��ȥ���F���u�5y+��=~[v�<�3���"���@3�5%[
�9n7?Q�������X���.���,��$�N����܆\]�����2x���u���MZ�f�^0�a���-��n(����'�%)���'ƍp͉Ͻ`�:��A�r$��V�KK�)��u9'gV�.PB\��.CvK
B�8l�ڿQ��PabtE;� ��1�E�ж+N n��|#ll���h`jo?��r�$1�*�Ǉ�^�z�?�H���P��W�fSa9U���klV�u:��b/�`����$Ff����镞L�.2o�lԶL^�aai�\���'�/er�!�[;Ǟ�_���6�
�.Uor<D|�-=�J���-��Ť0)�L)ȴ/��LQ���B1�Ȕ~XdP�M������xa�ɳ��m@'��(��x.c���O��+ć_��v�T7�i���+D�W�n�Ia������1�ׂ���+��
V��K�^T*|i&��G���+ᾂ��1d��ș��[�}�r����r���� _'���ϟ�V�g��)F����0$7�]�,`_dWrW1�Iu����2��ye�~1D�d`��
�<I�C�� /&��kx�����l� N��Ҝz�c�uUq�D�V�R!��'���{� jo��2g���sA�,R����	V
�K�h�"��'��-ϼ�V�k�Y�ە��p��dZG�'��ۊ�1zġ��f��:���R�,%��-�~\�=s�*v/�2g��-���<��~�D!��9����D�rμ�����z�%L51�ځ?dNXOf�cm�巬q�7AЈ4�fM��'?]Kd��>�8�u�t�چ�z/׼S�6G1V�Z%f�q��T3)Ԣ-��mW����>�cVJ���I a4h<dP[�7��sT������96WA����&Mw��w�_����.�=�bƚDy���l�~+O�x�#x�����%��l]����@��J�`{P 1��
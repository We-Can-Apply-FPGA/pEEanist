��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n7iE:Θ�u�>Rz����@x"�I�?���KmM�91�'0
}���Εs,NڍU��S:�������@ e���t"D%�7����>E]]0�j��lԜ�\�wp�\�W��@�e��^φn¦d;���s��Z�����XA�2�w9�E�I��Qx�F�A<�����c96O߻�w�%nƊ!B�����Vy�{]{��[�E�F�9�P�nj?.@y�3�{���s�RLc��?`��;�x1���.w*u�N�)n��L������1��Z������:�?��<���hw��l#�U�����@|�-�|�7Mg$JUa��F��l����{����-�7���s	ʮ%_r�J�u���s�oĵ/7�+	@	�\#2� ThiɃ������:���	|k]*���C�XFkv�Xx6�T��ȣ��D�F/i
v�8s��^l@y	�$��*��r�".3/�+���S���G�޶��Q�Ş2^S�D�����_P���F�(��~���s�M�S������A�j_懕EE�RB��+�����^�-"�t�t���(��+	�=w4o����&�4�p� I�$��KJ.|�7+��'=��i�B�ƈ�ء�/�c�<� �i���F����zkF���B4�(�@�i<�H���I�^/rT�h)���/��:'�n�.ه<��)�dAD�@/�z���^x]"l�pK�u��p�}q�eJ9��R�gSJ��5O�.�_��؄�w'1[�)+����L�;�u���+ ����0l�2��	6-SK;耷N�{r9�6L���`�1Y�x��_�%����]�c�d���L�X�wS�I����2�5J�z�v���w�-[���`
���9�)��}5�l�����{A�t���e^� j�#q�>zje҃-m:�����^��
�I&�w|�x�N�0ж:"k�Sf�P�� ;&���w����[w&���Ƴ����E5>��|��t\�BǞ���f �r��!��� hS�����7Δ������_�e�j���u�)�����$���p�`b'�e�fV�����}��g AM�)�9H��vq��!zO(c����#�2��4ΐ�(�i��v
�R�2p��
�D��&�:H|�NZ�	P%�e#cڋ����D��Z�i;"�2iH펼�4<'�� ���8yf�%��|!Xܱ����h�ms6�X7Me�w\���5y��� ,b�(�V��ZVif�_�"���#_E
?,B8���
�˭�%+c��!ܰ���4�׊�Y��Y��:�X��9��i�^ۼ2�V�O�<XN�T\=�{�fB��NS� a���=d�uW�N��������b�F�t�*}jm���B'��}��ͳY"EO ~�{r7�x��`X�_��ב+*���ê��$���9�FƘI&A?`�+�!��x��5V;���e��[I;��OBE*:=��'uCt3�p���lT�EZ�����OqF���7���]O�X����x�Q���OA���p��)�g�F]��O�x��<�B b\f%L6�,ε %� �S�#s��:o�ĩbp���wjy��?��9 TH�W��S��o3WJ�f��K��~^���C�8�$&t����^�'-�q����0*ya�Z\�zD��Ki�1>2W�}�T$����&p��+�����B�.t�X�z���/��.������s[�]1��W)%��6?� u%�,S���I4gu��k�<s�E^~��Y�I��%6�'���fT~����A�g��XĊr��)#L����v�q�G��<	~X�cp��4� ��R�D~�୾ĭ�>�B���3e+bܽ+��)Kc_�r�Z#Y���
,��B�6y���ݱ�MS���{]��;m<^���������f��NJK*��6p�_/7#��|�e	�re��:�"��.���� ��_lz<y�$d��3��r"���qC�Ұ�@��N.j��F�d.'p�ѳ#A'lQ
_�rv�jo6W	��6}&�^,v����0���,�+a}?u����[�Q��bzx�ݲ�yLd�YS��]G\���ս�Q��)A�6c�R��%�ϭ�Qq�~�3�����e�u�����~S��Uoڤ��7�@Y7��(nƮ2��TזZ�>��^:A��hkRv1�^����o��>��;�g2k��$K��y2~)���1���yT��ʎ�Mu�wa�oǒ�.[Q?��|�g�f�#;�Y!֗?Z�sg4.$W87�9b'ֵ'�:���N>K����J����	�&����;�C%c}������ �"���a�o#��t*��h�5�'F�i+yrV�ڊO��<�s��~$n����4` %�CdK���.Wd��G_�k��:�x$�a	�uԶ<d�5���ک;�jc�L��'8���
��ƀ�da��H���ğ����+&i�
�w7v��$�KNKv!�ٶ���
e�L���[���)T�tz3!X:�4�&"n�N�$=����E���f}����Q�|���0&!�g�ԓ���µ��D�-{�p��`N�dzg��I��Є��D�����Z��xz���V**��I?��6�lh�ٮ��_�����"pu�c������	03C�/뀗Q�[����&Ӧ���Y2�9iK��\_^o#J�����x<��w!Q�W7D�N��C·J�\�e_�ܷf90�o�S�(�p��G`��j��;�������ºW�9�S��u���'�\2�\����B�j��j���u8��hݏ�T�Ν$�~'�Bv�`�Io:�(�Q0M�!#�pL��#��q�0\�Z�+1�~'l[ѧ(�i017iY�0��a���Wr�W� �����%�:ӫ��.��\��m���}`W��|-������K�oC#Ϭ?%�}���;v��zT�;�K���ߡz�g0z?��K	�0���@�#�����Ƈ@���UD㿸@peΣ�?�V�YCQuMġqY�r{|�2+��uք	9K�h��1�$C��#h�����,��|��;y�wD�v%">�z�Z2������J����m�o+�<$���&72���.����k<v��ԉbq!�?��-5�}�[�}�`s���^+>$������hn�9�����^�"�q�/��v[3Ӯ�����an[lgu�5J���A���
�P|�8��e}c�3�53��ll�V��cB��ګ����g�'��!h��g� l2iB�/چSx�fb����ς:�����<Ǌ:À��%+P>�m�h��P�^IO])�����A1oB�������SCو:��}�F�o�E�N'�5Q��{�>9ya�G�Ι�"��
����'��2et�P�~-Fh��W�g0m��<C:��h�v���5�ӆgJ2��Z@���G�XnT����>W^Mg,ݥWU��z7`�����q�^�=-��˜ 5kT�㪴�a�D��5)��妨 A���������ȗ)�L[
-��zt�O�r$�vޢU����}�O��P���;�I�":Kل2#�'�Pt��	[�;�r	(�n��w͝2�ث�Gom�����р/�5�5&����
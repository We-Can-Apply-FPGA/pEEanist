// nios.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module nios (
		input  wire        clk_clk,          //       clk.clk
		output wire        clk_100k_clk,     //  clk_100k.clk
		output wire        clk_12m_clk,      //   clk_12m.clk
		input  wire [9:0]  fft_cnt_export,   //   fft_cnt.export
		input  wire [23:0] fft_img_export,   //   fft_img.export
		input  wire [23:0] fft_real_export,  //  fft_real.export
		input  wire        fft_start_export, // fft_start.export
		output wire        lcd_RS,           //       lcd.RS
		output wire        lcd_RW,           //          .RW
		inout  wire [7:0]  lcd_data,         //          .data
		output wire        lcd_E,            //          .E
		output wire [31:0] pc_export,        //        pc.export
		input  wire        reset_reset_n,    //     reset.reset_n
		input  wire        rs232_rxd,        //     rs232.rxd
		output wire        rs232_txd,        //          .txd
		input  wire        rs232_cts_n,      //          .cts_n
		output wire        rs232_rts_n,      //          .rts_n
		output wire [12:0] sdram_addr,       //     sdram.addr
		output wire [1:0]  sdram_ba,         //          .ba
		output wire        sdram_cas_n,      //          .cas_n
		output wire        sdram_cke,        //          .cke
		output wire        sdram_cs_n,       //          .cs_n
		inout  wire [31:0] sdram_dq,         //          .dq
		output wire [3:0]  sdram_dqm,        //          .dqm
		output wire        sdram_ras_n,      //          .ras_n
		output wire        sdram_we_n,       //          .we_n
		output wire        sdram_clk_clk,    // sdram_clk.clk
		inout  wire [15:0] sram_DQ,          //      sram.DQ
		output wire [19:0] sram_ADDR,        //          .ADDR
		output wire        sram_LB_N,        //          .LB_N
		output wire        sram_UB_N,        //          .UB_N
		output wire        sram_CE_N,        //          .CE_N
		output wire        sram_OE_N,        //          .OE_N
		output wire        sram_WE_N         //          .WE_N
	);

	wire         pll_c0_clk;                                             // pll:c0 -> [cpu:clk, fft_cnt:clk, fft_img:clk, fft_real:clk, fft_start:clk, irq_mapper:clk, jtag:clk, lcd:clk, mm_interconnect_0:pll_c0_clk, onchip_memory:clk, pio_output:clk, rs232:clk, rst_controller:clk, sdram:clk, sram:clk, timer:clk]
	wire  [31:0] cpu_data_master_readdata;                               // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                            // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                            // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [28:0] cpu_data_master_address;                                // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                             // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                   // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                          // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                  // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                              // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                        // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                     // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [28:0] cpu_instruction_master_address;                         // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                            // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                   // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;      // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;   // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;      // sram:readdata -> mm_interconnect_0:sram_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;       // mm_interconnect_0:sram_avalon_sram_slave_address -> sram:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;          // mm_interconnect_0:sram_avalon_sram_slave_read -> sram:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;    // mm_interconnect_0:sram_avalon_sram_slave_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid; // sram:readdatavalid -> mm_interconnect_0:sram_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;         // mm_interconnect_0:sram_avalon_sram_slave_write -> sram:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;     // mm_interconnect_0:sram_avalon_sram_slave_writedata -> sram:writedata
	wire   [7:0] mm_interconnect_0_lcd_control_slave_readdata;           // lcd:readdata -> mm_interconnect_0:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_control_slave_address;            // mm_interconnect_0:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_0_lcd_control_slave_read;               // mm_interconnect_0:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_0_lcd_control_slave_begintransfer;      // mm_interconnect_0:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_0_lcd_control_slave_write;              // mm_interconnect_0:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_0_lcd_control_slave_writedata;          // mm_interconnect_0:lcd_control_slave_writedata -> lcd:writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;         // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;      // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;      // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;          // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;             // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;       // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;            // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;        // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;               // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                   // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                  // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;              // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;          // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;            // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_s1_address;             // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;          // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;               // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;           // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;               // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_rs232_s1_chipselect;                  // mm_interconnect_0:rs232_s1_chipselect -> rs232:chipselect
	wire  [15:0] mm_interconnect_0_rs232_s1_readdata;                    // rs232:readdata -> mm_interconnect_0:rs232_s1_readdata
	wire   [2:0] mm_interconnect_0_rs232_s1_address;                     // mm_interconnect_0:rs232_s1_address -> rs232:address
	wire         mm_interconnect_0_rs232_s1_read;                        // mm_interconnect_0:rs232_s1_read -> rs232:read_n
	wire         mm_interconnect_0_rs232_s1_begintransfer;               // mm_interconnect_0:rs232_s1_begintransfer -> rs232:begintransfer
	wire         mm_interconnect_0_rs232_s1_write;                       // mm_interconnect_0:rs232_s1_write -> rs232:write_n
	wire  [15:0] mm_interconnect_0_rs232_s1_writedata;                   // mm_interconnect_0:rs232_s1_writedata -> rs232:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                  // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                    // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                     // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                       // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                   // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_pio_output_s1_chipselect;             // mm_interconnect_0:pio_output_s1_chipselect -> pio_output:chipselect
	wire  [31:0] mm_interconnect_0_pio_output_s1_readdata;               // pio_output:readdata -> mm_interconnect_0:pio_output_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_output_s1_address;                // mm_interconnect_0:pio_output_s1_address -> pio_output:address
	wire         mm_interconnect_0_pio_output_s1_write;                  // mm_interconnect_0:pio_output_s1_write -> pio_output:write_n
	wire  [31:0] mm_interconnect_0_pio_output_s1_writedata;              // mm_interconnect_0:pio_output_s1_writedata -> pio_output:writedata
	wire  [31:0] mm_interconnect_0_fft_real_s1_readdata;                 // fft_real:readdata -> mm_interconnect_0:fft_real_s1_readdata
	wire   [1:0] mm_interconnect_0_fft_real_s1_address;                  // mm_interconnect_0:fft_real_s1_address -> fft_real:address
	wire  [31:0] mm_interconnect_0_fft_img_s1_readdata;                  // fft_img:readdata -> mm_interconnect_0:fft_img_s1_readdata
	wire   [1:0] mm_interconnect_0_fft_img_s1_address;                   // mm_interconnect_0:fft_img_s1_address -> fft_img:address
	wire         mm_interconnect_0_fft_start_s1_chipselect;              // mm_interconnect_0:fft_start_s1_chipselect -> fft_start:chipselect
	wire  [31:0] mm_interconnect_0_fft_start_s1_readdata;                // fft_start:readdata -> mm_interconnect_0:fft_start_s1_readdata
	wire   [1:0] mm_interconnect_0_fft_start_s1_address;                 // mm_interconnect_0:fft_start_s1_address -> fft_start:address
	wire         mm_interconnect_0_fft_start_s1_write;                   // mm_interconnect_0:fft_start_s1_write -> fft_start:write_n
	wire  [31:0] mm_interconnect_0_fft_start_s1_writedata;               // mm_interconnect_0:fft_start_s1_writedata -> fft_start:writedata
	wire  [31:0] mm_interconnect_0_fft_cnt_s1_readdata;                  // fft_cnt:readdata -> mm_interconnect_0:fft_cnt_s1_readdata
	wire   [1:0] mm_interconnect_0_fft_cnt_s1_address;                   // mm_interconnect_0:fft_cnt_s1_address -> fft_cnt:address
	wire         irq_mapper_receiver0_irq;                               // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                               // rs232:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                               // timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                               // fft_start:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                            // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [cpu:reset_n, fft_cnt:reset_n, fft_img:reset_n, fft_real:reset_n, fft_start:reset_n, irq_mapper:reset, jtag:rst_n, lcd:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, pio_output:reset_n, rs232:reset_n, rst_translator:in_reset, sdram:reset_n, sram:reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                          // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	nios_cpu cpu (
		.clk                                 (pll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios_fft_cnt fft_cnt (
		.clk      (pll_c0_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_fft_cnt_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fft_cnt_s1_readdata), //                    .readdata
		.in_port  (fft_cnt_export)                         // external_connection.export
	);

	nios_fft_img fft_img (
		.clk      (pll_c0_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_fft_img_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fft_img_s1_readdata), //                    .readdata
		.in_port  (fft_img_export)                         // external_connection.export
	);

	nios_fft_img fft_real (
		.clk      (pll_c0_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_fft_real_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fft_real_s1_readdata), //                    .readdata
		.in_port  (fft_real_export)                         // external_connection.export
	);

	nios_fft_start fft_start (
		.clk        (pll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_fft_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fft_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fft_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fft_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fft_start_s1_readdata),   //                    .readdata
		.in_port    (fft_start_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                   //                 irq.irq
	);

	nios_jtag jtag (
		.clk            (pll_c0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios_lcd lcd (
		.reset_n       (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.clk           (pll_c0_clk),                                        //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_RS),                                            //      external.export
		.LCD_RW        (lcd_RW),                                            //              .export
		.LCD_data      (lcd_data),                                          //              .export
		.LCD_E         (lcd_E)                                              //              .export
	);

	nios_onchip_memory onchip_memory (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	nios_pio_output pio_output (
		.clk        (pll_c0_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_output_s1_readdata),   //                    .readdata
		.out_port   (pc_export)                                   // external_connection.export
	);

	nios_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                             //                    c1.clk
		.c2        (clk_12m_clk),                               //                    c2.clk
		.c3        (clk_100k_clk),                              //                    c3.clk
		.areset    (),                                          //        areset_conduit.export
		.locked    (),                                          //        locked_conduit.export
		.phasedone ()                                           //     phasedone_conduit.export
	);

	nios_rs232 rs232 (
		.clk           (pll_c0_clk),                               //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_rs232_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_rs232_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_rs232_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_rs232_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_rs232_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_rs232_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_rs232_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (rs232_rxd),                                // external_connection.export
		.txd           (rs232_txd),                                //                    .export
		.cts_n         (rs232_cts_n),                              //                    .export
		.rts_n         (rs232_rts_n),                              //                    .export
		.irq           (irq_mapper_receiver1_irq)                  //                 irq.irq
	);

	nios_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	nios_sram sram (
		.clk           (pll_c0_clk),                                             //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                              //                   .export
		.SRAM_LB_N     (sram_LB_N),                                              //                   .export
		.SRAM_UB_N     (sram_UB_N),                                              //                   .export
		.SRAM_CE_N     (sram_CE_N),                                              //                   .export
		.SRAM_OE_N     (sram_OE_N),                                              //                   .export
		.SRAM_WE_N     (sram_WE_N),                                              //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_timer timer (
		.clk        (pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                //                                       clk_0_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                             //                                          pll_c0.clk
		.cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                         //                 cpu_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                            //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                             //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                   //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                               //                                                .readdata
		.cpu_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                          //                                                .readdatavalid
		.cpu_data_master_write                                 (cpu_data_master_write),                                  //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                              //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                            //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                         //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                     //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                            //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                        //                                                .readdata
		.cpu_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                   //                                                .readdatavalid
		.cpu_debug_mem_slave_address                           (mm_interconnect_0_cpu_debug_mem_slave_address),          //                             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                             (mm_interconnect_0_cpu_debug_mem_slave_write),            //                                                .write
		.cpu_debug_mem_slave_read                              (mm_interconnect_0_cpu_debug_mem_slave_read),             //                                                .read
		.cpu_debug_mem_slave_readdata                          (mm_interconnect_0_cpu_debug_mem_slave_readdata),         //                                                .readdata
		.cpu_debug_mem_slave_writedata                         (mm_interconnect_0_cpu_debug_mem_slave_writedata),        //                                                .writedata
		.cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),       //                                                .byteenable
		.cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),      //                                                .waitrequest
		.cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),      //                                                .debugaccess
		.fft_cnt_s1_address                                    (mm_interconnect_0_fft_cnt_s1_address),                   //                                      fft_cnt_s1.address
		.fft_cnt_s1_readdata                                   (mm_interconnect_0_fft_cnt_s1_readdata),                  //                                                .readdata
		.fft_img_s1_address                                    (mm_interconnect_0_fft_img_s1_address),                   //                                      fft_img_s1.address
		.fft_img_s1_readdata                                   (mm_interconnect_0_fft_img_s1_readdata),                  //                                                .readdata
		.fft_real_s1_address                                   (mm_interconnect_0_fft_real_s1_address),                  //                                     fft_real_s1.address
		.fft_real_s1_readdata                                  (mm_interconnect_0_fft_real_s1_readdata),                 //                                                .readdata
		.fft_start_s1_address                                  (mm_interconnect_0_fft_start_s1_address),                 //                                    fft_start_s1.address
		.fft_start_s1_write                                    (mm_interconnect_0_fft_start_s1_write),                   //                                                .write
		.fft_start_s1_readdata                                 (mm_interconnect_0_fft_start_s1_readdata),                //                                                .readdata
		.fft_start_s1_writedata                                (mm_interconnect_0_fft_start_s1_writedata),               //                                                .writedata
		.fft_start_s1_chipselect                               (mm_interconnect_0_fft_start_s1_chipselect),              //                                                .chipselect
		.jtag_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_avalon_jtag_slave_address),       //                          jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_avalon_jtag_slave_write),         //                                                .write
		.jtag_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_avalon_jtag_slave_read),          //                                                .read
		.jtag_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),      //                                                .readdata
		.jtag_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),     //                                                .writedata
		.jtag_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),   //                                                .waitrequest
		.jtag_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),    //                                                .chipselect
		.lcd_control_slave_address                             (mm_interconnect_0_lcd_control_slave_address),            //                               lcd_control_slave.address
		.lcd_control_slave_write                               (mm_interconnect_0_lcd_control_slave_write),              //                                                .write
		.lcd_control_slave_read                                (mm_interconnect_0_lcd_control_slave_read),               //                                                .read
		.lcd_control_slave_readdata                            (mm_interconnect_0_lcd_control_slave_readdata),           //                                                .readdata
		.lcd_control_slave_writedata                           (mm_interconnect_0_lcd_control_slave_writedata),          //                                                .writedata
		.lcd_control_slave_begintransfer                       (mm_interconnect_0_lcd_control_slave_begintransfer),      //                                                .begintransfer
		.onchip_memory_s1_address                              (mm_interconnect_0_onchip_memory_s1_address),             //                                onchip_memory_s1.address
		.onchip_memory_s1_write                                (mm_interconnect_0_onchip_memory_s1_write),               //                                                .write
		.onchip_memory_s1_readdata                             (mm_interconnect_0_onchip_memory_s1_readdata),            //                                                .readdata
		.onchip_memory_s1_writedata                            (mm_interconnect_0_onchip_memory_s1_writedata),           //                                                .writedata
		.onchip_memory_s1_byteenable                           (mm_interconnect_0_onchip_memory_s1_byteenable),          //                                                .byteenable
		.onchip_memory_s1_chipselect                           (mm_interconnect_0_onchip_memory_s1_chipselect),          //                                                .chipselect
		.onchip_memory_s1_clken                                (mm_interconnect_0_onchip_memory_s1_clken),               //                                                .clken
		.pio_output_s1_address                                 (mm_interconnect_0_pio_output_s1_address),                //                                   pio_output_s1.address
		.pio_output_s1_write                                   (mm_interconnect_0_pio_output_s1_write),                  //                                                .write
		.pio_output_s1_readdata                                (mm_interconnect_0_pio_output_s1_readdata),               //                                                .readdata
		.pio_output_s1_writedata                               (mm_interconnect_0_pio_output_s1_writedata),              //                                                .writedata
		.pio_output_s1_chipselect                              (mm_interconnect_0_pio_output_s1_chipselect),             //                                                .chipselect
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                  //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                   //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),               //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),              //                                                .writedata
		.rs232_s1_address                                      (mm_interconnect_0_rs232_s1_address),                     //                                        rs232_s1.address
		.rs232_s1_write                                        (mm_interconnect_0_rs232_s1_write),                       //                                                .write
		.rs232_s1_read                                         (mm_interconnect_0_rs232_s1_read),                        //                                                .read
		.rs232_s1_readdata                                     (mm_interconnect_0_rs232_s1_readdata),                    //                                                .readdata
		.rs232_s1_writedata                                    (mm_interconnect_0_rs232_s1_writedata),                   //                                                .writedata
		.rs232_s1_begintransfer                                (mm_interconnect_0_rs232_s1_begintransfer),               //                                                .begintransfer
		.rs232_s1_chipselect                                   (mm_interconnect_0_rs232_s1_chipselect),                  //                                                .chipselect
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                     //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                       //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                        //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                    //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                   //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                  //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),               //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                 //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                  //                                                .chipselect
		.sram_avalon_sram_slave_address                        (mm_interconnect_0_sram_avalon_sram_slave_address),       //                          sram_avalon_sram_slave.address
		.sram_avalon_sram_slave_write                          (mm_interconnect_0_sram_avalon_sram_slave_write),         //                                                .write
		.sram_avalon_sram_slave_read                           (mm_interconnect_0_sram_avalon_sram_slave_read),          //                                                .read
		.sram_avalon_sram_slave_readdata                       (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                                                .readdata
		.sram_avalon_sram_slave_writedata                      (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                                                .writedata
		.sram_avalon_sram_slave_byteenable                     (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                                                .byteenable
		.sram_avalon_sram_slave_readdatavalid                  (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid), //                                                .readdatavalid
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                     //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                       //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                    //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                   //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect)                   //                                                .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

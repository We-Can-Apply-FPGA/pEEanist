
module easy (
	clk_clk,
	clk_100k_clk,
	clk_12m_clk,
	reset_reset_n,
	sdram_clk_clk);	

	input		clk_clk;
	output		clk_100k_clk;
	output		clk_12m_clk;
	input		reset_reset_n;
	output		sdram_clk_clk;
endmodule

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�8Ӝ��'���=�4m$M�# �2��ݦ"()��Y^�~���-Dѐŷ�f�b�����v�=����{�X6xB��Eh���ps)�s$�Ik>�;bVcs�r󕧱�cg��i9����@����=ݫ������q8���>R��I��Z�^��!e0�F->�eF�T�5%����,�
�x�Lz��H
q|���C����eX���̫N���u5�����Ҕ�]UE��$�����J%�t���BG�+��̊��;)�wcn��P�=��C�5T�7M �k���-��}���C�2``l?�ֻ#�:�����]8��m��� ��Uxy�r��O�b����r-l�+��v����m��! 2}U�w�q9�8�=���y��|#C:�������:���lNs�6M�l����6�t��Y���3��CZ�S����P�]�8�%�&�<��)K�|��f�Q#U;;�����I����E��A��rf~��n{sX�NT��5 ��fn7AHp�u���?6���uM5¶Y�kA����-s���ߨ�k�iQ�t�v�a��S�%�C�¥@��I�]��I.�T;�)ƾt;�E�~i^ܩt>>q��B[�i���0��`�f�ޑ���q�`���M�fRKo�6��7P�A�(q%��)n.��=���`��Mdc�d�R#��Y���-d���CKP>8�hx|��S����wq'�xopҌB�kz΃�Ȣ0J>g�8]uj`t<i.�m
w�H�&*k2$G�֫FP6�<����NA�Oҽћ�q��`Ľ�i�NO���vb����� �x����"Tt<��������uw���Xf�{�������ɡ�0#���1�7+4j�hI�Q�<ѕ��9�J�7�r�]"��[_/O_/��1{���-�?��P��L���K�����	����Q��/��P��1UU.��+�wZ��ބ	Թ��F*�6K�1!�%�KN��T����j]�jr���YY�<Hv��;;g?��� k�X������1�Z���	n�,gpNƑ�(�mW=2�u	ml렟��0RJ'ȯW?�Z��w�f^���&��S3H4_& �0b���6-�]��`ޘ��?Jb���>��cg���TGDZ5�.8��ͣ����qr�*��=c*,��q�[Z�ԟͳû��N�\(@��c����;k%���c���l��љb���r�B�L�:��lj�89=�8��$靯��rظD�7�?Z����{���m��<\���n5�{�x��ڗ��:+�;m�3C�@��w�r��`)�������)�2��f��c�$6��z3�
с-�v���R�Pȁ՜������N�tYm�}g�uZ��֚C&�g����{�4h��IU��/Ó |�R{�}o�p�I��Q�	8dJb`���HQ��|`���ك��qD��4b��FyJ����x��D�2:����b���FT�Q�y|pw `?�,�1�5	��m�/&�����ĦkX�����h�3�R�ft ����\a�Ol=mB��px@J�m2X���A� `�8�7cU�sqU�r��QJ�w���Z����:�s�ym�RahN��CxU��ִw(��U39J)M!��"*��): L�tY�D�d���&�*?P���ZN�\�v���KO��P+����[B�-�p7��,���h�;�ҕ�����|9��;d�Ze���Q*L��!ͮ|�>��ӡ"�p+)��h[�Q�|������=K^x*r5�����a�^7vP�6~�Pu�W�m��O�R�.@Km� �涳�Q�$��42��<)nh�e��M�� ���k�݃ǣ�JA`_��x⃼�So��r_��9'G�[���.�.
������y��ڡ�yM�M3��̽�|�-��>��~�ت$��p�A���923=��'�
~&�S���X�	�Nȇg��/f��*#g��6k�2� �uF'�2>�j[��h��^*c����I���CS��B/l��q�y^I��k���m�Y�[���D��M���ss����}���7}؁[N�d��R�qV4�j�/W��՜e�Lm�>��g�1�7!�Mf_��@)a�4x��I��kF��sI�,�c�g��� ᛩ���Z@%��lL^���n�L�A05�V����v<aHiz���N,0v���7��'�v�ܴ�d��$��Ƣz�(�O�D����FG�ILApmׅ��p]`?1����� (�����V�z�W� |�柹����̻��Z�ם(�µ%�[�р�h8·)-�Am�>�����H@UFA>�
���ںbi��}���3��~�mB�<�S����,b�y�Z�j�5�X�
���_���u�,���1�Z��*i4
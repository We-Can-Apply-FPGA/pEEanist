��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���nUbO��b��ؑnG��_�� �ݮ�J�d�o��4��ʌ��8�5�Lo�L",�,Q�A�NHc�$��|ฏ��w�f|�)lO/J�mM�/5�c�2Ŗ}�a��ޮ��M����A�d�hC�م^<�9�TkV�����:��)�x�ɮ�̼Z�j=�=u^�'�F�&k͹���Q����`�L�`/���v��-�������-��~����<�1|_��	��I�);�s�iV4���kn����_��:"�FN�l���1�48d[���ފ�ſ<̯���-�c�?���Z�	��F{�%�!^:���)�!Z{=*���d,��G&�F�f��5 5s�U7ٺ�p2�GK+R%ٖ�}<��!FX�h��~z7�X@<�
�tL��F4��h��}�'sHL�׾Qqk����$�Cq =�7�H�&�)��#�*�G$����v$KI�$YYSV�e`o�v�t��E�Y%��H��A��d *7�(���}��䗗<��̜KSHv�l�M�U%�֜4f�"p/�u�ާ��46� �g��!R�h �Drb#��jL����ս��˔ƢJ�y{UB����EBF�����bfD��ygD���`��i�yae�RK`j�D��7�$M����z۲�@����h6`=~������H���wAS`V�G�t��{�.���?��]taR���Bp!k�y���q�Y���m�Y�#w�]s�n���%��	��B1n0����u�Ѧ0��j�P�xZ��h&L>qw�zC
,hv0��e�:۩��6S��6?q����3��6m%i]�k����j��4�������_��Hj�ebSI�/����d2���)fLŬa��A����MI�8&T�jֳ6����Г����n�������7*<�JZ�}�,��3(4&N�릞�ΧQn�d��ڔ4�T�n�.v;���kK��..�D�mA�,�U�D�{����=k3�.��E~Gw��J����I^ci�Oϋ�<ۣ,$��RQN��3t��3簒�s�aA�s�&��!�%(Fn#KnDX|��i��X�hN�n�巚c��~�1	��ƈkd{�*��:�D�����`�0��=�}�����cH�gxA��ǝ�a�UA�;�	/Ų��jzz�qs3ΰ���$�9_�[�rڶ�u6;��pd��ގJ�K׸HS��ќi%�q�4܂�zRb]��2b��s�y��˓|�u:�>�L5ϝ��*/#;�7�6~�A9�|)l��w�ٍ4}���0��~�S^!%4�#��i_����\&;�	I��˞uk�q��a.�q����>�eA�>�-i!�K2k��EI.A�mQ����W0c_[���Pg�����R�K����7���/Ne�U<`J�ˌc�@JD�_-[�7
@�7��7�-f�_�)S�ˆ˙��G��Ю��b���Z��@f����.�;GǕ���Ҁ�Q�6 �u!��ߐ�0��f�Q�\�-����J(��{�J��mj5���Y��^-s�t섨���w�	��(�x��\A�i��Q���{�e�����p��(f�S������`�ZQr&�n�Ҵ��]C��)ǟ�]rG �F#y�����PC���D{��k��"����$+��@*�(I���������v�i�b�h�kd�(���#d����m�ϡ7��i����kl��$�O��Bg��33hv�_��kʂP����g��h��S�,Ť�98V]t��4�0�h|`�쁉e���htR��;Q]��b� r�e�5ז0ƙiT�4�[GW� lArNY��%����od(g�O���o�=\��B2�N��H5&������<T:��.*�v����A�����0�0Sa��~����uJQ%~i����ϖS\�l�����X��g�����E����*��M_�&x������p��� ��Zqz�����~�{�@	M���3Ѹ�=n���������s�s{�qQE�<�/�cHC��v\[D���Y�A�~³��G�#�1�4AJ�c����4��Ր_�dFг3�پO�j},�<��~GV�& �s�'ruX �|�=��gD`���{B	�Vi3v6?��ם��rM�U x�ϣF�gsn��!m=�W�D��;�X:a�&��x6�徺��M��`*�w�f�ج����퀲l�~�_E�l
%��ƭ��5A�B��^o���&|��B��)
h�;�X=ʈ��9?�������="�����D��U{���U�܅'��A�C�qW(�4���q��k�Y�yݼ�{oQ�ݓ��kDo������>���.��@��<��f�6 ��~]_�	�h�{�iׁ@lvͥ��]��zn�����5v(�S�/�'D����&)��P��Q����(������a3��+�@�:z7%�BR�&�ĈD��`��ֻ��`8�K��r2�(^����8`Pu��4���]��,��bE�W<��P�<XCՅS��,T�"�O�7(��ӆ������J�~#r�u�A���b��,��D~�晔���
+_;�LЯ����s�+�=b.ϝo*�ǘ@��ك�D猅&���v��v4���I�P�j&"K��yp]s��\)�Ci�8����]����α8$Q�YA���b֎q��	�d1�V\ʍ©�i��{��9L���]HKq�Q_O��v�����i��<��#�%fYZ����_O\��Y'��>��KR��@��Cq¸��"�ʒ��Y�j�_�9l�_�r��3=�����(�&���n�����1S��҄��:�Ub�ԥ�'%��v��ՂZ�|y<��߄���3}�x �[T6:�x6M�P^0����4�{K���#|P���2͸���Y��V�O�8�Sm'�c�:�U�w[��P�36�%d��	�U��d����p��Ď�(�q3���bs����kD����p?�	��[��%s����/�*�>�"|�0=q�X�(�ج��d���T0�P��9O8�,��-�U׾�[y^)��45���|�Շ���[n����6�� ��4�J����}�?�K�X��>��j��������A�X��]�F5�Y��*Uj��D���5�,�P����2��z̑*V�w�[�Au2(�U�,k;f򵷊~���-�3i��o����e���_=5��^��	�t�$����2?)X��N�ats�].�N�����Bث��[ֳ�����lF�v��Nk�
�:���Q)��n��U��Z�ejɂ�2o��>>�Yy�T���5�¬�7�iO����:��A�]"\rW���P�%թ���q$�PTYN�B[v������i�l�����Wǖsfm!�D��wIK�AWC�\n�QZ�q)�����h�O�?b�+<�&R�
`�}&�e6ᡜX¦�z#�Sdu�7:Bv�������\�j��[��3+�l�iAJ8關��;��TԤŒ��r�GE9�Q��^] �Uꅧú�9�b%���nr��m�-G3.Oj����;����L#8)�$ƫ2��:cGh;4ЭM|�A�`7e\�c|�l��{��^\k��YL��C�H��S�hTw$ ���s��	��>��KJs�J��6���=�x�_�S
r֘�(�w��,� ��YEH�ĥ��xi%�3T��X�"E�xsY�|Ԓ� �D��O���2�D��C"�V).�ί��񽘤9Vף'��Ksx�٫G��;�aW��j�O�=��>�I��b�n�o'\�aF�5e&IHƟ-���E�5f�V��_����{;�&0q�Z�4��-��ʶ�V(
���j�cS�b���K�����~H�Xµ@�����V������=b���{�i�y�P�Nk�X<��T�v�C��4U�2����y$�c�ۅ�����Gp������N��rYD7}M��=��a��\�<'��}d�t����8\#2��>D�y��=I/%�p��q�-�ۣ*���]���fm�_�s|����p�5.0C_�J�K�=_},*Q���u�yS̥�_�Y���m$���IN�T�F�EG(H��Xl���^�Oz�����2�����JL2�"5��c��MbD$���Ӄ�E:��ͪsj��hB�lC����f���sv�b�c�{H�O\��"������QŪ7~K=;��G�`�ǆ<Hx�G��8��̆��f`7SH�A��z�����/��:�Ľ�nX�·�?nB!�9&��$�g���ٙ�?�7��YE����/tG�l�(��>��P]q#I4������%g��QjV�q�u!�{��Rx�r�4��7�P���bs�%o�����{UFS|u���@�/�~�d־�-/aLgM*��l;(�E�]0�HA�\v���Ky�������m�o�'�}q��H
�<��FN����{��M����&�8Kʟ������WP�? �>��<N6���6&�>g�˞�y`��s�t1
)�U����a)��W����^���,ơ�X��T��*����5;��l�hAa,߷t�g	�Djd^$4'�3�B3�dD
~s�[)��3�@���4�f��=z�t�5E�*���S�.���
\딦�'L��8�8��:'Z#U�v))׎�'��A���g�.��.�t-��V����_�2*f���'�ʖ$C�Y�dd���Wqؘ�J$�_9���5*C��O�����:�b�P��34�hR/H.YZ�As����I�v������D�q����u�������U&����'-^u�TmqP�c��<Cl')�=���p�of��Y1�t�$�I�W��F���Q��g  &���!�/��Z�q/��tpD?���|���Z�g��0���]�h��|vO�x)%�)���7F�kδ-I�@~$��q�PI"P��HV�~��@�L��n��Ƅ��Ճݩ���wY�H�>�7��=ҷ�1�}�4z�Z�+6������f N��ߕ3������f��N�IjO����8���a��}�J�M,�{�=�Ħ@�LSp�Mv�VƮq��)��ITN�j�����Id�Uq ���U+U%��P:��r������4P+�}�#S�\[S
��z�H���i�+ќ�5�ڣ��ukd�?�ܛ5��(�Z#
a�5;�P!��=r@Cg2�Q�d�q.�6)���hJ�ai���*����T�4o���	W��eYlKo�ܲ����OWT�G���U�+��=�mx%H�O��.q%��)��뀁Q��+M�)�����N������>�T\��]��S���{������[\X����+����}d��.2�*SSv)}�)Z��AT��.@�)KDI�<z�h�ֶ�^�_}Νnc���8j�̅r^
���Y�H�v�+Y@\�ln�jw}����ɓ�Q��>�
�p=�Շ᭶��N�Z���4�?�1~��'A�:�=����S������ct?��mɒ��2�9ư��حް��Q�1T)S��~!�
o<yHI�ƭ�i8Fx;��wd��?���s�	��%I��i�cap�Qʴ���6�_%����@��+�N��ʈ�@�֜��l+`�����k�<���&, �ӏz'op��j7� �x�,���CT;��9��p[7�^�� �8�9��D�>Հ�;���Ϩ-��U$��v��@�,|�Y����8Ž��z�;�� c�"@Gu�l�M �����~;6��--yW�I�1�܆���R�t�TGky�3�I��1&�v-�%'t/2�\���A#Hf��yZS�2��v �͎5�ݿ�J>��7���wt�J����V�|�?�X���̱��=e5�� ���-��T�ZZ.#�F�� ��2�}C!MO��6M�����͇FHƋ*K��O�;��r `(�zݸ���g�kS*:O.K��fnLQ����H@��s������M�L\	pK^J�$ d|,��[]�J��^T�����o�J�O��)��������
Z���L�վ���D��5z���qn�bֆ�B�X=�5�N���d�C�T��H��[<��va�����vM���ŋ�M���G�d	Q�s[
01�~�i�H�M�)�/�p�*�^�s��1)�^�_CG�
�Z�1�Ѭ�pj��5Zۍ�f�h�вqE��wEZ�L���0̑a	�>-�]e�r����p��K��Lx��W�Ъ�On���j�ɪ��v@�Tkѹ�����MT?�[gKZ�������&t�&%��O��4��<��})Ű��!.�q
���t��]*�4!L0V��}βD�&��bO�;,�V�$���N2eֻ}CG{��$�9�t��y�/��q��E�!5���6��؅C6H���@�^ǌ��7�(���I�ҫ�d����B��W�s4��uH�{��:5��CX�r*V��rZإ�X;�������nUT\�G�����L0�^�G�n;�QSE���6�����k����E��L޷�a'�_�+;2k�J{.��]��Ea��T1��U�z�ќ���A��݁1�,Jc:?�\%%��+�y5"D�d�/M����>F~+�q�X��Vs���kM'�
�/~�+��n�kT΀�������QZ�*�|�k�Ut�YT����O 6�-�M�xws��vGි���-$U.�M�Ȗ��3*� ��Z�wL����a&ܺz�ƣ_X�]��� 1�����`�濚��4���+���ru�J�ؽn:;'j��q�.�݌��*�Ěj�?�"m�4�\g��  �1�Nצ�v�ĝ�i*��(q9XE֋��\�-AA�ܨUZ4���F�
9 ��н+"�&,ث����y�Ɓ���Fb��&jY�Iz�tz\)�#��
=k�ߛdw=O���'��Ǧ�w��h�hʨ}ݷ�H=M[w�Dc�Xc��zǂ�[�.v��I�`eF����F)	i+UwT���·Wc�v�~��Vn��m�<J�p��G�����]����o7�}.�%x�@�����J@��t�f8���*�d�I���]�r��,���a�pꢃ
 ��FҶs�?KJE����Ne�?��۷�9���#�M�o]��i��?PU֭���S�$��l8~���t�C�CJ�F�R�P��P�j%^k�x�N�v9����E/AQ�Ͳ�תS/�V?N��b���Io	Z����9�U*j��l�������v��YP�Q���9?��1RW�XhD��:�>4�5�e�Wz =� ��I�g��!@�-�Up�z���������p���ex��?�|�0ӌ���z��Z̖ ?���QE�0�c��Hd�V�w�
mG����bAS|�iȻ8Z�6;�]o�H�e����\�eqzBdmrӃ8��,R^��Dz��P~󛀔��yA. +S�w�9X�����@�1�g�4��P����B��a��&�)��u������Fn��"���5��we/���o5��"5(>g�\_�Tgr���'U3�"�mJ���X;����J\��r���-�b�� �|ϙO��q�u<m)vB���m�ȹz*�4��'�Fb���h@�����u��[�A�ez,އǻ��b流���-��
����۹���/t��Ο���Y?��n��u�~-�u@3����er���b{�6�`�*��� ��9�֜�Y���PK)(0�c�W���#[u�$M���S�4�"
��R��z=i��З��oem-	MY)&��9���:�0��3h�ɂ�
��:��JM��,'��@���>�9t�h�UH���P�\(���N\���ږَ�gS�!��4�]!��H�^P���T���\Y�w���3x�F�.�Ņ��Y,0$y��E���k��]�<�b0	b���j(6ܶ�lL�:�}���Ƒ������/\>�����%\�tHj����֬���)��B�y2�u������WM����*r�-��+�_�ģ�0-o#��(�qo	�8"a9h>q�d3�����G�y�y���No�����)�1����x�3���K��3ME:p�v���*��t��+�+v�B$2�}-��l�'\K�i���
����#�U��5���y	
�￱г/����ZL݋;:nk|�+>�l�`	�w zN���MZ���Gg��D��O@�T}��F*��53~�鏈~�ÿ��=�%�Q<4���ͨ�P����&�t�ioXAm##���/�H��;�˶�2��q�y���,%0���l��	��L�O�тQLv��$M��-_��Y��s��ؘ;̢T��s9�>b�~�Զ^o�?�&{�U��T��w�\
�UVY��`����'x_���o����x-��ZW4ۏ�Y%,e�ٙZs���9�*~F�����O���	��0C�a
D|�E�U����l�("�b�ba ��\�"�V^Fx���VP��>[�KHB�8kb+0�Ի�7�\_���������
�x,��d���A5��P����7�4��(6�<�H8	8\7�����lV~*p�.�.L��>�m�j5 O������,-\K�}�ӽ�L���	��2T�yY��G�EmYɋV!�FT�,e�)�rS�	����ռ����ĵ�<u��.6�W������Ҹ�J�#ZY��ꭜS,�#y�T뺖��a�1z��j�+���K�4��[��쀠"�b�?�h���VZ�gT��Zոu�@���7+͠�n@���F>ȬV�Pfv�Rq
�=�O�Rw �ȾW<ܨ]����C��hWERt���9#j�c�Uy|�&�b��d[6Ǳ `��	n��m���F�V������K��ZKSl�|N����Un�;�[7�5Hߒ��a�-�WP∣��U`l�4��k��9AZ�Y&�F�-H��=�$�[)��{��k.[�p�x����h��D�������#\�움�~3�	���]���eS��S�xb^"�A�����EX�bu1�k!��iB|m�X�vSXb���W��R�10 �+���Jyb��?�[+S�Xp�=���\�u��).�/A�3a�u,g?TЁ�~$���< ����o��z[���r|���T-[�S�@��풉�λ���аDIj�B{9R�B��^�:�G��	xƊƕ"{�����dZz�9�H͓k��)R�GL������-Q$��!9nm�\��o��i��3�����3�^%ۼ����s��1��V��g;��fi�?��O|��}�����+A(�T0��Z���ᏪW�Lx�W '�����3�jN-�dg��9�-"�j.aV�C��U��q\�G\HHV'?�M�p�R.���W�_��:��Uv����	=�2�Ps9e[S�ܡ z�2\#Sb_�B��SA�-���>61^������w8C3y����PD=�� Tf�G�qh<s_���jG[�"U�S䫍�����F-������E}�����˔8�L���t�sM~�)ϙ�u�U$Έ$�j
��~~2�����"eZ6�kF@ c�+�h��ǎQ�ثPd�i���mM�u�\� Y\pWNi��	R9�/��J�!m�v�~��Bz�,�Cqf�K���BW�x��`�Q��'L>�Q髆�+47�\���T�a����^@�VZ}<_������g�\�khϋK���g�t���g(�,̃Ϥ�<.�R 4�7s8Z.���^u�ez�Ÿ:U1��IQ�y\bʵ��QS:h�k�-%��y1?���E5�mC�H� �i!9I2œ�N�"��0�E�h���; �s�p���r�$�~��F���@��l��ǐ�1;�糂s!���A�3���G�+�=�/1�Ӫ�T�K�ˌWA\�v�2߬FF���3����kp�X8�;�Ǘ\��BK�3A�y$(��OAC�b)����x�(�!�C1��Na��g�46
̳ u��n^��B��}��Air�5�ߋ�f���<M�k������1�,8��� I6��o��[qᨌi}cw�L��)Y�#�Gj����ڬE�N��`�wY�T��p���U4]T�!$g�m��<7?���U.\��H�m�O͗��V2�Uwn+�>�ʍ>���-L�W%l*������] ��w;�!�h���0�wFٰ�lw��>����;��uNc\.����Lc3j�,�m�2b�kR��|~��M�m�t^�w����v�7 G��oH���x"l��L�fu3�KCy������'^���E�VV����2��������:Qw������k�B3)�(��^��� ��f��T@�0VD�9����ý��,{3�}p�� -[=�����?�c~��z��~�f��;	x/����r1�#|��u��Hj�P�{�RT1ήwu/H$X���E����C�����d�0���#�d&� $0�O�A?�1�iMdq����F�(���	������:�p�όgb`s�(ԫ ZI+_:��.�Y�C��M�'�BX4�N�Q#��uZsz��e!?��!�r��t�P�L�ǷԞ���$�ޗ;*AlӨp)�ˢJ���T�P��ۅaK����A�$�ï�cxY`}#~B�)`��;>� Vȸ��T���~���u� ���UT����-��\���%F�i>L����,f��!i���"Q�TpU@j�FL���sbP���jB �?���d��������Ǒ���=��#�k�"3ҔKFO�3�7����iѺ�t���7�bS�"�{G1>�-�9C	�ŋ��p�V���U�׼���3����*�ܿ�)�VE�s��[BV�X�'�U�k��e_��BW��g �a����*\�ϞSdiT�"".)g��'��|1z▏�9Ќ�d��{F!���%Suv�0뾽���b�t9���`��Ae��5��}Y�O�L��<w�)����B�2YH�
|��M���[r��8��%<n^���a�J}RTt.����8$d�v��ζ:;��x��V�����b��﨣:�"�K�xv�r���rg��{�!Gщ��]ֈoۥ����d�Lr�}Ju������#ݨ�3x|�@��;╧t�Rc�g��߂x��64Fn�@��.��G3��jmdv2׊��j�Q�`�h��Ԧ7��(���E������P9zsl�e���ô'<'�M�V���)�7�B�����a�8�"�2���ի�?:
@��b����0�r�l���M6�M�azc��x��Kc�{��,�+C\���28���a��ڶ��ե���g��Ln�maR��	W_C����]�_)V{��	�I��R��a�mȴ��*E�#�B5����E�8�\JCF*���[��fn�����)Wi��7�C�:6�y���ރ��~�탉�;n���2�Rk���t`Yߜ2�L�V9[�_�A&Ձ�z�� b7��H�m��|��<0;
;�6��?J�q�9\/C�q�]RX��J���y?DD�3JgeX���1f�'���#� Z�xgÖ���e{�U3xd��^�G>а��'?0]��7�0�GY�����X��Ra�Db�������DQ�P%�5M���H/9�%�f,�� �Uy�a��v��3��4mK� <����P^_㦴ě�+�bD�9�Y�ם���i(�ѫ6>�I�fq�����]��4y�ug<U�.����0���>�͵�L�\(���c�W�H#�,E�a���vh�X��0S�1�kJI�ɾI��^��Fu�u����z�?s'N(��aR>g���R��[�mѧ)hZ1�����5ݣ�zU��Z�����M��h?�)�[��z؂�"���zp	�S{]p������}�&i��#=�[�7�A�X$=�� ��_$��gk�M��f���N�k��QYE��L�{��p5G��'[�,��?���O��F���%e�ҩ�;�f������|��l��K>���9��0�h������Mg���j�i�������J�Fq��'�"I���삱��6�Q�w�uS���s��UtK�T �'&�
��� ���_�7[3�Xb�@@"�jh��/�偝Jc��}5����W�c�w�Z+3EG�f˖���D6@j]��y9�#����:��)�:�1�}�2<"�tf�gn�ʕx�w��
�4+���]��x�k
��E�$��mq�k�Q���vO�;�i���0��B��;��.�C]>by�S��,0_��Q�� _����p'����D|Q/8[Pd�!3��$xT���5���k�o ��:���$��=A���a+"�m[��� \xW:�jú��/�&�똖�k�����(aE=�'iŲ�G��P����WTA7�$�6�� F�m'�M�!��ٵ��!����4�<C����t=I'�����čXn#z�n�J�՛��[S���^����5ޠ�݉e���!��/�U1�M�r��I����7�;''���W-���w0a:AQA�I/`4�U�܉V�3��hB��Ŕ�\5�0��К�(�Ω����9V�Dԗ���,�T��v:x@��=F��ږ���M:B� I[�?���� �p��z~b�@�G��{��ݩF����fk�}�ڶ4��@SJ�=�!�b�T���o�1e
ceQ��x��l��8a�9�#5Yx�&��mO3�Z@\��W���Ml>�Ϣ����ǧ|�N^[�	��k�%��������C��~�H���f��Cƿ�q��傰���j��9��S\޲�o-s\�"����i/9.�)m:��lDspX����
�:�.�k�X�)����|�Ų�u�R�� ��k��P���E��{ �� ?�,�)�r�i>e^�v��z)|�B�bŎU�L�6T_ie1��}����a��F8������q����x��0a���j ��π�����"�9���
c�� ��	��B��B֍e�l�H�s�����}n�A�{��Uʶ�)�������C�t1`HB��B���y�'��R ��s�m�,u�J�j���'��P�������$�l�w�T=��~��BJ�D�m$׼s��	���* 	;j�$
�����;�ҋIе��Ow�_���P^�RD�&�̸R���Mi�/E�1�kH��Z���7hD(�k(l$���r�3#AK V�@E(�Q��U�Йn��s���6c��J`p����+2V笫�,�
W��O�d{:��%�^��'ѳ�|�G����ڭ�G�K߱qmj(A���/�Ojw��� ��-qf�4�Z]����WX%/�V<�w�f�e+���jm�=��A�W�3B��$���1.��P�/��u�,x�+�ir=���s�� ?
�e�w��s��%�em���l�����ih��g3�D���1�r�Fx)�6��������&����bP0f�ـǑ�Β��>���	�`,�TBY7VR���?�g���Q�x����ݨD��`�p�I�0�{�����:��x�����֔[��k�^+���:BC2\{�>�a{�1Rp���J��?��ĸ�Y���k��(3}\�S.E�(�-�Ov���������<����/�@,��.R�E�0�CC�߾�n�B/J���g��?#�����0��)f
���fnU<���6`W��9�Nt7�dd$�]J|������ �l>�������� Af��xOv����Y�L�����AIl��f�%@���� ��� d��[�NԨ�R0j:B���!l(�|F�WơJ���J�����3˫#k4z��~�l� ��%�Z]���H/1c�[e�(�R1+��r������:�@���������Ȼ�n����{Sl-aW*'���, ��:�����bb�"�]���	<�F D���>kb�(>`�4�s�ǖ{�0�K~wF\�P��5�f�yH�"Pb����	䙬*�,�� ���h��0��0f�7'� u.�L���nW����{���a�+�u�J�7a��q��S7�ђn�s����6B������;�C����M5	B��C�$jx��]����!��݇ܯ�[_;A�K�z�>��Y��bU��CI
2V�ݲI搈{�/�����a�iu�.N]q��-�+ ױ�{�<��0rqdy�W#���f�Ⱥ�yI��Cbl�>6�̚�7�O܋����jd(O�3�v�(�2����5苏%�X�����4���6d��2��~����v\����d4�N�����_�{����D���.�QH��(�&���d[�g�F>����ә�S�k]����@!�.��/'�9��Ƽ
y��_��d� /X@�_q�w���r�Me:���KH�Į]N8�`gR}�ۈ{8'$S�Cx�iTc��|h�4V�z�>�9�W��w�p�g� �޴ц ����D|�u��J3f,�-iy�˵^@daڤU;*�E0ܣSC;�j��cU����zpT�L���_�>9�&Y��M[9�<=䈒qV_��D��]�	_+�O�[���<���%/��m6�@cOƘX��7��xR/L뎣 47Q�v�{'GX�ny�	#C0��p�1=܂�.���T$��AǛ�a֒J�Ϲ~�f�r*)}\;��>@�k��C��O�� }�P֢5�j�bDb�����k'e��Rȹ����{I��Su׿���r���9E��/���9�®'�_>S�"�~W(�D5�)�C6r����ފZ{.i����n�t�"<�c�=³"��+t/P�~�X��d���ãu	��
|����dz�R<nf����X��y�,�'~���;��g�KS���ߍ!�������K����<�T��@�Ji���^ϲg�?qI���G�tm��{2:�'�^��t]�e�O 3U��Ld�q1l7��rR�j�e�pD~�R�Vɐu�7<Y� B����)�1��wA��N�Ȉ�m3wg*��S�����1/����ca���Z�A1,s"�a��`��s'�C/Pk�ϖ0���B�,�.��ZZ��u�5�,
U�$g-��o��Vy�J�"+�J��[F(ej�_��y�V�_��)���QΘL\�������{��0Gc ܳJ�8���0pDO�]W�����ӟD]���O����I1�T�r~��d���q��~ޟ�4���١���
���ЊD��]�8/s ���E��w� ��{f~ř,�WR�WU��)N'`��C�N�8���*��o�{�g8��o�O�f�/KOH�۳&M���#�Un7�3�v����5��V۠�h#��K���)M��,�i]�V���%���\�ލ�O��M��/�ؽ��.�N�M�9��u]#(� ��`_�<�z"%�j�͊��k��:5q=�N{���ײ ť��J*��G '��3�ؼ�Ep�
~&}K��.b��T�^��N����Эzq���ʕGb
�uYL��"�y+Ч��2����_�̭�f��fՎW���EYZ�2d���9�R(*$���G�S�E����[m6��3�@_�P�9 �jh��Ga�bW��:�׽�90ԟ��t����Hn�C=����$eag&Ќb(D'�vD�[��o8�b��tI�\$��
�P��3�"�*��A��iX Si;��9�yq���d�����g�*���
 o;d/�9n�
�v�YϘ( �d�\op�EU��ޖi��>����u����u�O�+�9K�� N���_�_��픯��2��5E��h�DF�F�tfDmw}�%�
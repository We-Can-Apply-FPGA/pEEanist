��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i��������쀞L̓"�oܜf�~�5@�g4�5�	�
����,aeH>)�3+,���KԾ�D�X��x���ark��!��H�ҫC��\���!Q{���,�1C��g'u��:��55��$��%.�3 &�S��EL�V�a˳yUҋ��)�33iG}�ɶ��*�'�_Tɮ� �������3@8�B16�@�
����_���.����ʑx�]�_!&'�;Bxl�a�Ɗь�B:�b"��1�R-������TbZ2qDT��Ԑ�2���d����]1"���-Q�ˉ��{�03D%��T�H:N�-ʔ�r|2K��}�T��8n/��TX��Y��fB��X��#1�7�t���D��_J9!��1�B"��V��Q�)��Pi���D�s)�2\�~�I_֥3�|���hv������t�A �7��x��1�� ���״�s
~�*-d�hu�֝5?���eL�L�.�����f�1�T6�.�ɵ�߼>�J�
�
b��%9`AЀ@�x�i�v�J�6�W�L_#�zat�B��-�@L4}��߹��D!�F�S8��k㬪ґgK��R��5Z'�����֒A�0"��V?�S�v�+�˹��f��)�]d��q��1'��04��n�b1q-����g�����F.)I�E�|kl�î�t���>혠=�;$<?���A��{�j���B�X�\fpEC�U-�7��?DX_���uj�Ⱦ����ױ$E`40�Y>�
^C䔴��#�)-��j�������H�\��=E��jZ��;Tϒj�b<g%L�����+) XQPĦF[���4�@Dg��QZ#���6H
ǽ�2͖ �_/o/G�ɦQ�*�]}X�Ϗ���m��=?��u_%	rB��������^b͛�����ώ]93���BM3_��s��f�e �Aĥ1G�㮹����xJ�H����z�p�U�*1�\.S�K�Y��{����nq�-i��L�9CZx��]3�*��Fd=Z������#@g#��ש����
�-D�Z~�?��i��}�%����n��1�r>�B3]��}���	E��i�\��tg�3��-1V�b��� ���~�}�%P��L ���܊~v�1�W�n���l\�6wSDMYYq����vP%� �)��C�z=G9��-����z��耪����'����J#DxY`4��0�z�����cq��[l6����}�\�wSFӵU�!v���'����m���*����&���]�uݗ��EQ4���x���x[�L��� ;�|B=���5���q� J��g  62:�8G�Y���S�i���K�~�v�.�㪌�Q����	L�|�K��緈��i�*�J	̒C��*4[�8�A�,ͅ���6¯{�#ةGԵ}�g|f�@��CY0���>���}YFskE������<�s�W{�ٱ��dF�i���E��Dw����_:#��#�X�����(��-8�����k�v&� �nޝ����S��N����*��;Uӓ)���P�Zc�g��w�6��OmM�Cz�q�!|�������� M[rݎ'c뙔�>�,!��W�͐rF�:���RT�%�Aʇ]{��5J���)c�`�{\3v��Ń�� ��@����L��Wff��|[4�v�y�]ܭ�j�8� �����eN���}�����@ZH��;�t`���E������uU�5����O�<�	�U���baMI��Q=�8յ��^��+�/ӊ��K��%w>���<.�A���ʺRE���Z_�x�
ͣ�7�P���!�~���tx�H���ju�G!Y�-�KX>�8��*�:w��|�o��o�J=h6_�6.�	�*\A_b}�m��T�!���=PX��p�ߥd0�'��d� ����Q1yB������p���v\��Rx�_�w�ԯX� ����z�$������aȷ�����l�|'����tw�.,���)L� 9g�;�EO�Q
�\���2M0S�ZQԆ~`wCB��!D4��	��5��en�|�^x�R��o����3������֛<��+�-��-ߪ�n�&����G}�F���B��nǝ^�'
S�û�=���d��T)[��b�/Z�"�
/�[���#u@A`���#��7�5�~�>'J�J��=�!���=5�2������޷ڟ�$�7{G�����rx3Tt����K��Ɲٹ���Y��5�"8Ȋ+��u[L$�\�¯'�Q�= 
��+F�'jϩ��_>XV�����S�w�o��v <�|�}3���M�<h*�*�F��~��Ωe��[�I��#u�?�<:��Gϯ\�)e���Xr<V�$(���`��`YAXĥ`�ل���> Ib�G�#�8�h�U�ʧ N%0Ŧ�%�>���e�8/+�[�����G��){���^�����05�y�3s ��د�I���J�/,<k���_�X�+���~F|S^��ߜ�=�N�I|��罟AJ�2Ƌ����_��*ԛ#T��mΥ����m�������_�.X�g>Ό��Z�x�":2�;�7�g'$�O��Z�e��Af��弸���I�y�0�}@:����j�z��~�οN����P�a�V����O�P\
�e�G�������H���ߜ�*�<Z��4�un5�����%f0O���z���Wp%��#ݭ��."��4M�J��fo� 8���O���� (���7Gq�����O�)�\(9��5]:��Ȁ®�Ky��b�����Jץ��Խ���!�Q���!q1OZV��Y�߀�dl���Qֶ��[F�Y�gTJ~��Ǳꐴ��K8��g�>,��r�i�D��X�^u:8�G��]��O"D��p������ �D/��:C/�O}�<ݸ��1:��W��U��͢�����s�%?)��֋,��<��������Ġ����>�snmr�DG�'����S����5���>{�>�l����mT����gx���=\�D�.ړ 	��Ģʚ������2�A�ZI�.��A�x'�i�p(b���͢l�e��o���vL?A�L���.=\xr�Z+%l��>f�5�oyf�V��2*Hy�A�{�*��:��5\н^��r�k�v��I��%}�.�?��:�nr���`w�Vy� ��JG"�+�$�3u��㫫�Ǵ~�J5�ޖ�S~e��k�'�E��#���4:;Y�b��Q`���{�!�D��ZF;�6,r��S82;t7
��f���*�q}��[~L���-�&8�~R�QW��6%~�}'u���[�ݬo2E�9������l�o:𭚏��J�p>��^��b#\M�[5+
��֒��I�Ps��Z�g�d�{B���o��C����k�]���k���Z6��T$���YB��h�'}=!)���C�A��BfKr&ӂjY����o���-�Ie��&q�B�/n��B����%"Eg�w�#Ş�C�c���وx��۞ϒ���4��'�)��m%_Q�۸�_*+z.�4Z�A�$Z��h��ɽT�(=�����	�I�6N��u���2�zw�����'��_�]�u��l>uz�7Yn�$m�v�5n����l�J;Ӿ���ʒf�u�_���UH��:í?`�R(����;��5yF��ALAo���N�X5;��0v�	��Wi�N�6�K���c�gJQ��!;�*�?_4�0���c�Aw]��4�w����jn[94��а����)�?�3��"y�j( S?�*r��d�K؋�*�TY���&��Ka�W�Iy�}=>���D>q���b�G%�Y�=Tն@5��Ȱ�tp�m�J'?����F[���	���]��Bv:E\օ	�b�7N&ȭ8�=��o�d���F/ض��u)�d����c���kW�e�f)�Y��A(�5�W����U]���.���cfy�JA�jI�ɓq��W�T˧�����������v�A��L��K�6��cBn�0R��hm���*	�Ϸ����m����7�k=>u}=r�J�&A�t�2��'&�n.1)0�hx�Q��F�+���aw�j*�D ��=`�h�E��;GQ*���V6�S�������O�.���M
�N�:(�UUiІ[ٯ��$QF�2�Z�$���Q'rL$챿��X���9L_U���}��߯�Y7�-�YF߅����_ڡ�'�� S�j|���ODs�m�9�o��5�e�
d���޵�
+��u,#!&텣\�b��*�U�w_ܝ�l�����ѧgT��>a�\��o�*���,�v�g�׆Vu!a˟*��G��#A`hA-��M��e�	����/�T	5S�s.����X���o~�7m�^���LP�m�c��z�5��Jr���{ 2�g��>�1M�7�)�?���'�]��]B�당i�Dϊ\b����F��5m�˰�4�8Aa�(�~�{^]�6R��+u�Z��A �Pʎ�А�\7��njh��7A�^SA@ֽw���q�ߡ�ٯ>�,�s�֦��� 0�6Q�Ui�^��Di�Fd��rnZP\��E�'\ G����������}��G���A�~��v�a�祡^�7�u}�
�[h�+0Y��l���X�6��*z���`�T%@�^���(v��Q=_��x�%Ї3��32).QS9-ފ7K�}�q"o��uG�E�;�N;��C-��;0e��s�-n�It���?Ng䧭���R��;� �,#FY[<�\Q��(	��H8d��(CTu;�����[���8��-޻ٿ�x6�h+��m��@ �~X�6<��d�(J id������SA����7�\�O��תi�c�ñ8�f��1<@��x�]��^V�>6��ʇ%�_��'����9�1��a��_��d�<�ZH֊g�z�}�A��C�x�Ͷ���n',��v���"��_ӈf� �{6 �TpG�$�1���	���+F�=�f�Ьߩ���ŗ�d5�s�l�(ry���@�h
T�J<a2XN38uHC�]%�X��� 7���ɘE��?Y��Ӏfp�
�"���9yL|��Ƕ�dE�8p����m��N��
�l�h����E���`�^U��R ^�L�v�~��Xx�p�b�ø}��!�m��O�-ْ��J� ���G�چ����Gj��׈����#��O
���Զ�j�\�d5���v���H^�V YY�e��r����X�Ȟ�����z�@�.X�Lpܸя.U���'�JB�l�xKT���H��T2HJ�p�$e0\*EC�=�!$1�7s�!����r����A�mg�Kw�����?��4�i���6s�7dx�������Qc��� rL�1,��0㶫U�b6=x��Y��@;��?b�[o޽�+m�9��/�[����#<�c�U�*lC;�j�3�I"x�	z����wh��&�C+�L����@��?��cd<�w�zN�$��+u��}�G���/��A6��q1��s �BZ�wF��Tc���=�
gO?E7�"/�F� "V}D���Ft��3��b�OL��b=l�I���W�%O�R�B��o��g��������w>������vr�h���Yyz�n�Wo4�n��jB�e2z�}Vஊ�o�J8��f�@ĺ~���9��^Օ"s�[/!$���J�/~��mF����Y 8������p0�J��G�k��X/SA����y[e;�&���J�8FY1�eCN������Ih~-��%�kA?XLО��dZ< 359���>�G#��],�0+�y���p}C����>D��7���RӦ~��Rb�P�\ L��'��4�6���������q�mpf}�_&!��ְv����a��+񠶂/ο��ж/|�~�Q�~���ZoO�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�
#�i�MS��Q�
<B
�t?{�^�z����$�����Yp�Z	��O@�/iO۸�3�����p�`��#���+�B�&��Tf�O�}�li��x������2��c$����<Ԡ'��Hb&�[�q8غAC
f������8��]vʝu����@���-@�0{o>����;��9���1!(�g���?�
C9
e�Y�[� y���Ts���b��Qu
�;τMk9'i�=���h���\='��c��+����墍�n:<��UN0��k��<j�[�ȋ#+a�ݨ���Y�z�cc�PK�2�g��yt�)��)�,��r[ú�� �_Zt-gpzR���֐a;c�պZR˞{F�kr�*�,"�e&P�+;7����]|�P����Ȳ軦��*�P��o��C��l�ب>��o���i�v�wMXq���s}̐(��}�c���MrLMʃ2mr�����t̄[��s�@��ČS�f:{|7{�,H���U���b�(�K��w�[j*��j&�=��Q+�n��gދe�(`0��$�A���w\��^7[AGI�TF�3�nZ�Q���e0�?�u��_GS���1�FBKp���P(�U<�隘�a(*�@�S�~M�3(P@�0큒`���F�X,��^ۘ�2�F
���9�(ol~�/J�(�f;�
[Ż���[��8W�실,�L�Aj�"x��ZY������8j�^�E[�]��`c��F��:���N"�M��Eö:5d�ul��g�{y�M�j������}5skX�Ɍ�9�oșÓ��f�=*�1����H�N�1�eˆI���
Q��8�1��댇2�+�e�
EZ�k.�J7��/��QwzwYt׵{�����x�p+"vc�!� l���pJ�:bu7��N|� +�Ƈ8i�J(~C6RF��
.�7:e�+�}�o���6�%(�������sB�R��43�C(��0�e�0�6a����yY2RZ��NZ0��i?�����H_\-�������fy�l1���jW�$�sp�n&�~��s�H�B �B�8�ݪ�\�vK����r!����XA��ڼ�g�r��
�L;;@Y���m��S�z緎If�������i;�k�ݐ����3�]����)�y� �ʥh�j!Ԓ���>�9Ex���u{X�h�dDE!�9�˰!��:�&��&�P���>�E�vQX]g[Ξ4T�ݡ`�3�?��~yW���XQ�n�W�d�so����r�Ux��e���ҧA�2y��0>?������L�p M����� ��b��hݤ�Գf�@W+���}l{��;1ʧ��r ������++���b���9��򼉃t���>���PYG��`I'�X��W=ةr��9iSKE���&�#�WhP�5�x$D��ۘ����)����&�-4�k�5�j�\�j��T`�Fݘr,�+��ы��L� �lG�Rl�T{�<G��|�]m� v<�a߲��%�X�Rx�\��M"��f';6	@�5�]/��n+]�0�E��)��r2���y[{��en}�<рE��f��V��w�H�}jh2Ve�c�(���;'in��7�]	)uQ򯿿�.20)m8h�`�а�Jbr�=��y�M3�3���<�o,A�oG>�I>M�
 4��l�b`��t����e= ڕ{�;^�ߛ�o�?�hI��.�Ы�<���8�{m�ZM	>���Ǔ?RE�A�a`.��S�[\
��4lp�xߟ;�F�p��[�9XzW�?k��V\1���4ϕU�	#VGU�tk�"N�빍�w��(��O�į�F��}��T�h��U@(�)�-�B�H
�a�%��I���<N���9���b^�
�,�E���_ڒ�w�%xA�2�~5~en�b��S��t��߭��� ���3,�.uB���T�r�u�u��vx�����Pxuw�6w0�Z��B�'�I�3�Si�A�Jy�l�W]�-]͠�t�ǋy��G�L����]*��4ҫ@Y'��!�[m	�o]~�u$�~�i�Ɋ�����d��z�/��� ���5�yDV-�q��=(�ғ�z�	��k*��\�M���Y��W�ɤ==CE#���J&�Wz�J�	Ԯt3��!�ĀQvP�8��O���64�GS��?�V�	���N�-$��i\�+ܽ��]��j`�T����ɛny�s�����Ǫބ"h��'e�x����^q�-���3ҷ(�$8�Z&�����7t �� �?/��p'�XZ��L`y!�8��d�c��ի����B5R8|��~oy����y9�q���0Ƴ�moz�Goa^�z�߷�613����z|yn��&�<���Nry+۸���.��7��'�iC�Ry������]|�&�iluo^w�ar�QjT	��jvA'pJ�0��r'�E���8%�c2���`�>"Lۡ��^��?,�ǄϠ&	��ʬ�S�������3`y�%��Vmd�={�(�$,�FU�-`W}�]�\���M'9�fjgRD��l7O'�,�0�� u^�k�s��}Q�:'��?�YU�&uд�.�:���&�}���}F�f�7R9�9�r���y�DN�|��Ț��{�|4��*��ʺ��kG3�TW�!�*C�����߸���Uω#.r:�"4���O�&�9�by�$j��^�7rH�g׮/���1%`�Y�wei��`<5>"F`?͜M4��	1���A����R~��:æ����VWC9�>C���\�ES��3�����ۃK��
��p܋�{78~�O�M�ytδ���͍����Rv&����N��f��䅿"�TYш����,��LJv u�0�5��Rd���hb?X�8=�ӓ��yr	�2�j����՚<��A0�t�����7ޘ��P^I"�`��f�����G��K�[�[�u�)	P�����g���(#��O�*0�*菁��k�n
�B*�#A�����(��O:��TP�J�:�<�`��x����0�zl�0Cw�;��N���5wc	�2�֘QV^��Ւ�"N��-�Y�1�@��f�ҏ�
)�,b��Ԥ�R!�d!#
�� ��m�F���lk�Gm�f��������S�]";��K. �^�2�n����D�*��)w�f�߃$j����k:e�*�λ�L��7�	�Ⱦ)��EoJ��C���;:��̓\�� ]�
C(d=�5JO�2���^).�FC�3*��۟ɯ�7X��.%��t��B$:�D�0RM����p<�!"�g�>�����1x*.���u󫫄����{�tU
Vw�:A����[�D�Q�Lpb��q�A[N�G�`N�_d8*�r�:�P`y�J�>����fi�=�7ZK�Ê坛͚9S�ӹW�iQ�eڨ�;(�b��z�L�qv�rO0�qķ�������c���ϰ�xNg�>����ҟ
\�� �爞���\[[��ɵ��|�诱o��x�.�� (\��˔O��P� �/�*D�����]�E����^�7�[���0��K�
�
��-�o7�B�-�Z!\�ѱw���&S���ԥN�UeK
`P�ϳ�~X�O�%��s6�?���%�L�7����ح���}?͑�k���O�>��mɫ0�z�$zWj��r*D�ڹ�;9���R��V$#y�����a�h�@\A�r��ML�`�ٵl��]꒠b�ʺu��/	�em��f�i�	2��nØ�Z<�X�N:t@��a�$}�Q��u��Gf-%�i��*X`M� Ϧlf~SHIn�q&�%�{��y��BJWY�(�X~ R��5K�_��$�C�>i���#�˰�2-6�ä���k��i����6��}�՛��Ƈ�Y�옵�����C����{B+[̓�� �</�h�W eqb}��џ���\�[Vd�I0�=d�`�&���p�n��&d=��v�"A����k�Y���Kn�U��D��}�������|{] �mZW�䜑ů;��xPL��p���̙܋2����LB։L`��G�?�+#^P�Y����� fI��~
wu���~�����E�M<��4Zɰ˚���+\5s�MUW�,�zz�:oxQ���VL�b,�}ܐ.���(V����G����{
���%^gx�2>�SōwR� ������3��a"r�����	��cE�Vf5�uj��*�o���t�ZjEz�����IL��'x#H�x��H��� �T�E�|B����&�k���J;�j۞Y�L[�X�vn�ɩ��A(�D�ܪ�h��D7`&�?�=��Z��8&�]^֞�&���DG���@�q�����S�Rv�n�5�IIRt�W���ȼ���=�ș�Y�f5���DKZ++�ԫ��\W�,�[q���y%S�.���P۴�ZFo)��4K`/*,@�O툼v, �!�8����6#i�NbZp��}�Z����jk�+Hy��~��  �Ë1(��w^A��������D�__�H)�
V�ޝ�
�7�2���P�L��vyr� \C���I�҂���v< cA,�v�I��7��ó"d*�]L�!���a;Z.��;�����t���@�,��Vg1�!�AE��й~��<����\����x�sҤ]�g�jc��@�V���;���fB?b�cK��s��!�ޒ�xhD�Q�Բ�qS��@��NŁ_0��2��x�y)�P���i5NP��Dk�gg���xGh�@$fqCk�+�i[Ӵ�o{q������s��Hjc�:"S�o��8q�~\���2v�'�Ž�[�]�8�P'��F/͐�͖#z�K��Q>�x�����cS(��J4���˃i�1�FN4�M�(N�Z��M'�6���g֣���z�?/ �>H£�#+}��5���7+
\
�T�B﨡i��\�i�J�OC ����J֥�&RF��m�Z�ao��@��X����9�A5�,v#���kє���b��ZP��얣B��QN"@F�p�WżG-��%�u���SΦ�R'���l)�m�ݺ%���0�W"w�*/P��b#��������ʐ��!3��%O,��R���~X^7m�o	>�!���)���a�4?w\C4�C���E^`��Q�"R���?b�h:�/�7��v��>��J����r0�7��w���R�b�~ʸ@��]�2c�cV����։C�`��ڋ��у�H\�^-����/���ں�cȪ�bs�/X����Er2Ѱ�+'ZE�K�*;V�ܨ��As܋�A��J"l�6�������:�>f���_���wgԦ����:�l.\��b<� ����
'����秔�̠�%�c������w����\�M���F[�=i��d�G��P]�*xY-�X��o�ypC����۸5j�A���q	�B�)�C��������@aR�{.9���>,���.#�
�B�{���B�+ψY0<�n����-�r��%���j�JitP٧Wk�VW��!6@_߲�5���8�J��ƍJy�7�$����*�T�Јx�Y;����Z�d�W�2e��f������wE�s�Į@���qg�^Au�/s�ډ���lF�����n*�K8�����hmb�1m߀�_#l���(XǶ���5�,���k��2\p �J�N�� ��&x�f�}�Ҿ�;Ef�O�:1�
/ͭ	GR����`�bѣ�H��`V�	�х�_��楤���z�ܹ�|z��˒�P;�1A}�g�� �]�r�]�ɞ� �-����z���4Gj{�&04��S$�d�'���,�z;�*@�#nK
�5�,�s�Px���`؁�*�M�l�Z��Y����Jmss��(���'��Ͳ�=a��&KT�	����;��(7��8KT�\���* �4�a��hfσ[%?���v�'��#�S�s .ݷ\u)�&'��G~P��%�lW�e��Vd�]��[�x���a/=����K6<T���b���<�\r*�����33d
g�mc���V�~#�8X�3*��|��L�OX������������9j*밮���� }�˽��.�÷b�f�L�MI���Å�-8f�/,���[�����Sy�z�R�C�h�w��1]��$N�r�L�h��B��~�2�~~JN�3����M������>s��H�DYהl�ͽ�����e����D����C��h�d�
���Y�'����N�a�M17��!��E�x�xe�3:ڡ��Ͼ"�)����/y�c��ˎ>+�O��	D�-J�j���a�px&�{�a��]ǂ�l����P�W==��HhH���4лx�"��%e��j�b�v(�� �}.�Q}Y0&��x#=�$J9���^��~;c��D���=Tv:����D��y�c���I�quz���B���`Gذ�P��'fBRE�'���#�D�:�e����s
��[z��p�M���J���b����z~�HL&=�[�])�u>`@3^4�,D�e4&��l��b(�ʂv����EH�{;���v�6���~	I�ܴ[����-\V���`����������6'z�r�ظ!�P ���5;���~__r_���~�9�8�P�Gp
*4M�R[��,����f4�fHD�w�yހͮx ��Y�u|�{%����Rs0)
��;
���u �_*�6O!�|�̵FϴɆ-������[UC��p�ЙWt~&����惞�Ѧ�"�'��1��a�����"�6�4/i'`Թ�6y9�I�U��@� -�
@-�B�Ź�W}jė�#�V�\�H�H �z��(�a�Ȭ�@��o�l���$���ܪPuA;��ԮX
yṛ`�o7t�A�u�?	�	Y�6D����P��
|&��k��'�C
�}A�hIfs�i�^r3[���9y�1Q�oW��Shr��P��-#=�M�-���@Uij����=Ůo3��ܛO���P���l��t:f�f*�կ�����1�أ��󇶝�&��P��nH�tKL������YfŢO��+m�p��
�~Ӊ��=�c��%�35[���G��.���vS)9�ą�<y1CPiL�@�)2㨻�8�9bhN����P����m_�X�9Vh�<�b���|������m�y=T���a�|�h��$��PN~�l{�����|y,S▤�;3k:mL<@��b�ų��n}5����/9�GI��Z�s�B��Z�@�,OvL���Td5$�I�M�l�	s���1��M*�X7����C/Hw �������L�rDKA��m��P/��fw	�F��ܞ'Q���5͈7t�&��c����~0�T�yQ�X������eɍ܋R�����w\A3i>�K�p��w[Xuzy^���"��`��G�?�W1?�D����	�;���j]��v��u�6>[K�[����\Xeeg{\������xȭ���H٦��V��Ke{s���@��y6f�wN
So2���Ĳ�c�Z�]��i���-6���e�0�ZSz�v�DT]�r{�Ղi0��(���"1������\J�^w���0�E�@k0���S�!37P�I�K.��)^���TI�	��:�f�S�-�������������4*E8��6�ܩB�-��Ps���/�q��-�y�W�s���nW��F(�Q<tH}�������&̘ʏ�
~�SV�����z>SN_#�	�8A�� ߚ�{iR�B��/�2s���V��X!X���=���1�Ι�ڲ4�C��Z�"ī{j޶��$��%A�I�ćZ��u߹�D�}8q�*��@ڶ�@�==nۿˮ��Cס"pWx�M��Kqө��K`�Q2f�s{g��
͵x�Kw
\�üch���;�!��[�r���+מ���	p�GmR�G^�g�"_��D1yփ���DD�̧��F���̀�D�fio/�#]<����c&�Z��f�����(�B-��J;&�]�m<=�l�G
����+jN��kJ�JZ�����!8���/��ɸh���Wq�z!CZ_ �}97O�A�]03�����y>��fBC>ȹ���`�|c���zZE��˄R��m%���m9�l=%i��tn��Tn�ggi���p�z�`�,ӳ��Ƅ}s�عIk̂�@�\��؁���z������D{,]��BY���8y�O)JX!��*��Jj&ķd/����8Ր�q�-�ko������'���������2�V�>>qu,�ʇ�螸��)�bw�M��) ��
&swXq���+�@i\��l(��E��
ׄ�-��Ƌ����6�2�LB��<	WU4�"�jl��ZnS���d���v�xSEyo��<�+p�=O�+��e�\���`����}Ip]������L�b4�7�����|�p	�`�(
��v\N<��ù�/GΏ��ci��z2r�OZt[<z��0�4�8P}�����XSmjrC~jl*�UI�R$���:�`�#ȭ��1�+�EX4-��WyT��pN&]'^Ƅ����ѡ
R�u��Ƚ��-��<Y�#x]�{˘t)���D�����b�)�[��~y�*/)Ħ��B9�B�.��S(��T�S�����n��q��愎�ߕ�![x|�f�&mV�9m��ðW�R�/^�}�Du���q�?��zP�^�W��k����ҷt�� t�)��K�9�`F�mA|W@;�H?	
"+�C֒z�[����m�M��3瘌�"�\v�x�H�U�{�����M�����f��Gd�5�Ӛ�����|����sm%${�Hlʂ4��S�|��GeXI0Ⱦ\�WZ�J�����?����l*M(-q�lE�GMX"��c�N�U=!��z1����hO��'�GZy��QK��Δv�Ϻ	�wM_1���4����c���y��~�2(��̓w��$U�������*'��$�$�@�+V�Ou�{3�HW��K/)-` ����E@v:�>\�6a����=َ��ԝ�RX�b��c����N�O�tf&smYK�}
d�B��3'��{�;Mi�Z뱵�S���
d^��\�,&��Xb�Tg�}JX %D嚺���뺋p�� ]{g3��ek��&��G� d��J=��|&�m8;�G˺��8⚕�Oa��-V�E3��k&���_ȂmN\w��\�Z����X��gyR��u�����j���������n:��b{`�i1��w#Wf�~Ƀ_���������RW�H:���>r	�D�V��}d������,�Z��2�l�R�rH��������l�88.9�A�v S�.��w#��
�v��z_:�3�A?t����M	��B�@ڲ��4�u ���HP���8P5�5h�Ɨ�(U�w�+�����2d��"������u�#7!�Ч�l��R}0��k1�N��d*d�~�T�ulY0`�0Ο�$hۨb��-ţ��=@׷%$}+3�6�fvW-Fco�\�V���Ե �����t�ȭ�Wxw�|�κ��Q� ��G#-5�7��Hi���u�(�W��[/y��L�#��t�M��s�'�'��e�4�K*��n�X~��Hت��Y�]��!�o϶�!��y����ŘX\���OUQ8h��2fL�r���d~VH[Y��l>
]��4�����{�O�ql�x�>0�0��r|F�O�CM�to���^���.���B;�t>�DOj����y�t�ΐ���,s�x�2z
zB�W�o��I�KB̥Q/����e!`ǯEא�+!h���ۂ[<'��+.�mB��m��y9)3h���*�,?͇9E��#1�M%t|�����Y��a��.�
��d�������t>H��!�T9 ���-\��
�'^)R����������*�R$~<�q���&���P��rmf���y[�s����*]�S���O�"Y��d�n)L/�Cǩ��*ճ���`��M�ؽ���t^�Hͱ�DMqpys�DW������U��-���é����s�nڭ��~|���uy_�.��1/�U$rI��L�j�H`�K���mQyƂ��={%{f�#;������k��B��T�:�	dV��4��+^��&uc�8���"�=��]R]�'���Ց9.������c%�9P!�N�$��n�eWɱ�GOɎ
Q P��1��^�z �)�Y[�ԜÀ��;����r@/��e���`׫d����K@1Sn`��c?�0� �$�F�<�_���[?CO�I�U��3RUn�Iu�j�/�2+���O�?���-���h�Zi�2F�H��<�{J��jF�<­�r�T�kV��М�2��<�$̭��	\��~��]q�d=!5�%�/ɖӱy���l(�Y�tc��	�'�0H$�*��l6��d��^>b�~��-��S�։�7�C*�v*�NN�|*�3~�F��Ɨ҅�S'���*��hŽ�h.��=>5�JK��[���6s|�C�a9
�5��4�4���@ݸ�Khy!w����D�೘�g+���?A��ܟ\��?3աe�s��B�r\�$�r��R:��
�M���*#��R�
L��ې,�+��v]'=x���L1l�os֎]�=C����G�$8�Ϧ�۷|,/�bGg�g띹ԳO^�_��ԯߠd*wi@F�5�:,%z��0�h�B1sS�J;����Ō��ш7�S[t���:�"������=H����0�C����p���g�P7˫�f"�f��QX��B�e@�a�zY��bf�5|3~������Ŕl��,�u1+��
A��9�8�0� �ׅ��q��98>$~�5����~���t���$q��.:h*p�3n�����ҽ��L&@�֓���*dt@�ܓ���9���:���6��>�dRYF�����t���sL}lW?������9����sdh�R���XJ-���N��N]:�lx��i����h��fMZ�DB�;�
P�>����sr����x6�t8��;���f�n��Θ� HSg[����� 4��NX�_�$�����N !
�D�`�\`Of~pJ��|�'*8uY�9���?����)0��û�^R�fz�դ����/:�ϸ��J��P��`u#2.�ͳдc��_��m�#�Gr�������c���{o�9L$��䷁f^���,�+���X��.Y�Ȁu}�4j�p��8���	Z؂���Xw쌐�E}�����2�%�E2|��z�3VK8[�sxJ�EA�2���2x��ۈ����fq�k,�aG�C]�V���K���V-|��*��p�@Z�ʗ�n*�}�D@���~�g'a��D��!��D;?��d���D�_M��x��j���8���n����8b��Ȑ�
omr�5�/E;X��������=(�2�R"�y�V�s�GSK���2�0��g;t)'4	mnl���b~�T.#�����fA��1�~a7�Qog�Y�Ri�8�4C���j�:�y?U~5�̔��g���E�3+�5��mC�iF`��I�Yз<t3�/���.ԣ'����4��AGdѳ��+`��r�Jj�1�I=�?��d��ʋ�\ZĎZo63�Z~c�w��+��1r�8#[�΅�t��T/�)�}h0H��@��G,/Ƃ��~R�1˧�Ƴ���B�@���o�@o?��� ��Y �1e{p����<�&@A�B3a] o�/��x(�Ǫ8�/kO���WmPޫ��e�r��$:��t���H��[��X�*xM�ջ:���au)��0ی����,mt���_R�L\�]b��ٱ�<Ŭ��Bَ�FU��L}K蛨W�0�_��D/ �lf��QZ
�e���pI(Θ�G���Kym[��_d|PUFӒ�r���װ��~��_*�k@�n2#Z�k�1K���ÚBz&�P��P�.�e�٭ʺhD��^5<���dM?�v2MП�-�����:~���+#̄�{r�#�@��&f<{��<ejױg"n;����+-�-�0D���R����5��<�6֕fn��(���|��RGg_��~�vٵ�s��@�x�]�KԈ���ՅDk�Kݏ���t���LL�P�%�TT�n�k ,��K��e4}xer2Ϫ�A!���V�u�i▎�,z���5n+�S�0���e���^2�VC�m��<���@�@�����$�-��.Z�����s�A�9��iXe�_lag��l 6Z�|`����)t�_�g� �,9��*N%SRԊ}s�*׋(���c���T�h_u��,'���h��$�d�����\�<�Hnϋ�eB�i��w�YU�������-�nUNe[G!�j#sC���Xь�j�:��Ǩ�[(���#@i��n&hr�F���s�A�t5���3��X�p��KGX�`���T�.��!�Jٰ``
�'A�,�]��J}���q����O��U}�mM�]��'Y�\���i�S%'�m�V��zYx��E�n�p����(�Zj�
����8�Ǫ��Vx�n�C,�R]ϼ_��/Ū,�/�΋�8�������ƾb��b�BTE%��w�\k� )�<TSnǋWc����V���d�
b\U��So����Rd&�E8�3�GF��{f�w�|����"�8�<���?(Yெ���B$^?c�3LƳy��x���A�i�V.	�G�c�`����a|���b�B��Y�O.¬�j����e�����-�C��#��V1]�n�#1�(]y��"���=��q,�\��9F�V�l_~/:�= h�҆�!`Y4�gP��&�>�u�B�}-�ǋ(u��V������ oȍ����t���O2TX5��z���� �^���;Ƥ���G��F�2�����p��m3z;����zwѷ	������	�^��wFB��׍�ܒ�fqy����h�Ϛ)����t|R�1��H��_g�s���|$�伇�&��Ѫ�J�B�� U�w����NhӠ�<���ܵ����1Ż�� ��ب�i� !!I��|�n+���e Ɩ��>����r�1�����Б��f��S��B3�D���'�.d�F�������X�G&\}@R�R��W�
�m���/sD�aTb]��f/�pV�p�� w�~��~l@��b4&/�6�0��*�(�6�0-l+�)F��8��崨Hͥ���Mۼ����%����i#���4��O�%1:\~� H���&�A������}ł���H@g�Ȇ~�����1��DŃl��䉐�+S���dP餱A�A�?8�5�/��3��7��bW�~^	ſ�ᆃ�D��\f).�4�t2�8��">�z�?�_�y�>bbJЇ��d��DR�%n�l8`(Vha\�����S�Pt �	<A�E21���i��~�˱X�霏�`��}�I|�����/lR�<9�1�@�ij�l�m\x�(F�R��A��O�=�ňۮ�:�ߝ��L�&szz�;Y*���`%�r$���j� aҀ<i���p�/4s��W{0JiT��2�W4*�Wd��7����W��0��h����k�`Oҧ}�S�a�?�:̋J��;
O�WU(��1�TA�6�נ��6�F��v-��� C�,��#�K�P-s.R7�)���>|b߿1�Dp\2���|pʉ|('L�}p���Q���l���K�����6�F�=��z�y���Oe�aHޖʢ�"���M�w(��Ж�=����S�rݝ�{P��S5�]�Ɔ�K�=GR?�J,�L�������9uM�x3L���	�+?X��c���l�Hޗ�a���w�G�r��]l$<��-�I)k�i�S�&D�����ڇZ鸵v�Q�6�iی�8r>�~���	-#ߐΏ��:r��O?�֬�������3�XQӾ�v6\I��ًߵ�{��Mj~$$��<8m�����~�
�d��J	��I��6=�Q"��/�'��F���鶰K��s2��,ퟔ �P�������q2����@9g].3�E��:J��o�?�%.l�_��U0���<t�m�-����2b��Lc�+��)W�5��A���hP֬O!'tk�"�F���,Q���8U>��y�K�doG>��,g1NW��&F���cR��썻\�H��C)f�e'�_t������������bh:aG��;�Q�7AYGy,��q� }v�X�>��f)��MFC�0U9om���.��Gn���Z�������]��xɞ�O&�\���pSߘ	�����	��uV��D�2"9��"8�0<6��ַ���#�5F���D�f��q�/�-�����}A�^�:r���1	/�R�p�ljֹ�׻*�B���V"�/��u��0�����M�Ix%Yz�"�ك�`�ƍ�-Z��4��Q��W1���G��ؔ
8e�Ľ�u5R��0_�"Mx_�9����Ũ,�S��y��猹M�=La���?F��a�cL߫��!��	 3��������8n��'fo��|� �����#*q���0�{����/�
䝁��ȸQ������';/o��l�Y���f�Rx��*+�C�u���J}m���Q5:Z��B������qV���d��2�S�� ��^G����i��G�C�C0��Фy���;&��-CM��k5��K�?�=��i1�sb<���8^sZi�@K���x��/�l��C�F����敼�<�e����P�����{Ti����.#��	bm0H��fB��mL~�R[Q"�6N6ݒ��	#�/gs W��]4�
\�c�v�I{O�/%�2�dow+����X�ua`����h�L�(���Y�J���%�Q2�$PQ!1��f������pØZ����w8-#�E[�ds��2~>�Xh����%�E�)���t`�����ػ��
�[����UuQ��蝉*��,�D�<_~ya	ؔDlf��ޔaF˼F�?uK���
?9�{�z<Z�di�R�y��2Y��~v��hD��1�4�'� �x�"]�ǈ���Rn�ՑU���}*y��OP��>�弚��E��!�?�q�����v�܍�n���@:��m��}U�XR�3�F82y�Iu�Y�&k�K�����_dK>��YW�B��;�YP���ζ���F���d�fbJҵ���̄��տ��oג�[7����G۶�s���f1�H��<����t`
�"�u�����W� n�)���aޮ�8@!���0	�-�/�҇)/��9�/�]��	꜑�K��vn�݀b��d���`Bv���� M?�ɵe�D}|���u������@`�J��{cÈч��3x)����g��D;�j��n�R���&,3�rB_C4�`scU�M���*���a�����>�pFaWP��$����i��a�����8�y����w�@N\��o�z歮����#2��q�N����ӛ��,t>螖��`�k2�.lFv�C�g(8��Fc��YݬK���G��|&v��ͳa6�h��@,�Fʂ�/�_i]^.�s��+��PO_�B�'QK��r�%�(�0�-���.)���e�'�FP�����t�E����uj����`�;`�3�?�N���xv�~�gW\�����ǖ��_�����y�EA��D������$�X/����:�P��j���ײ3h��"�m�Ã�*J���D��ܭԲ�����W:"�3ᱏ�j�x1�Z��O�WVA<<c2�'���B��6�A��-ƙ�X��4����ĺt�+W+0�#�c��^�ru�s4ک���z �t�䭶Srז8Q�sF����g:J�����I9���l2�L�T�(K�h�s�-�8��J�L�.n����KmV�I����Y8Ԏ���hr?�ך���yps9�-˺�7]VZ?�0�ܜ���d��g|�����݃K��&��o2��󸡣�j��1���܈��LrOc�.��~���+���)o�i #eF�G�����+g����wJj�`o�kJ�ތ��I8x�b)O�g�W�٨�X�Wp�ָ�?�d�:�qn��
�,6g��lB�'���]J�T�516-�����h�\��g�������,�C	4�R=7~q6i�5�ʥE��]֙�|�I��zN6�UPF����L	��8tL(f�v��o�L�%�4A����-x�4ܒ�Xi��I��6��g��S�'��j�5kc��WG~�^H���w%��ʥ�JtlU
O��6�_�6���	�8�.!���@w�b˛�����߰Jn0�kh����!�_�=�ǁ`y�'C�@/�.e�B�d�3NZkJ��ݴ�՘:A�a7��ҿ؏�̛�ʢh���SL��[��R�
��	��jS���B ���g���8u77b�ޑ֤%o5*3hp��ʍz�K��4�'靣�d��Vf�>lŘ)E�y�+Ի��w 9F{b)M��js�q(\3 �&�I�-1�����!Mq�������v��8`�)�mxOt���^�J��:�+S�n=���=.��U����k����;�n8h�������Y�^CG\�[����/<Bݐѩ��3@H�	�7����R�n�R�D`�`�^̠�������y�T�;>���5��2ӹD�`��O�ׅc�ȯ?�fm��ːn��m���/ց��	�����D�ú	.�O9,��'F�& �I���KS�
e�qo�B� � wc��(�[.hW�B��=����V���q��W�o�J娰�,#�ws*�K)��"��hI�-�ᕣ��BC�.��iR�(*$���e}o��p�榢�.8� 6�w�!͟v0�( r�!1[,�_,�k�VumU��3N�����
ͷᒖR���7�<��� d�봈52���}�*ڡ��a�W�k�lT�)���O��|����1��0�jD$�����^k͑�è���O��k�ؔ��b� ŋ�c���r =9n�ag�&f�Ƹ����N���i������$�����pg[��5�7x�t�ֶ�Pu�蘾�.�br�W�O�(�N�+��7�+�3� �Q�dzfNj��lu��{@Qf�3F�8���:���u`��d,� F"�|��o�n�Gr�j���vf`ǰ/�6���F�9��Ù_RaO�r+�N�5��Ӓӳ�du�|>��2��x�<V�Ϛ=��V��U3�^ݯ�c�la�_�����l�}9h�@�����;#KKV)���d�n�A�}��r�n�C�b9�D��=�A-���t&IJDZ�����1����!������+|���Pf-�ٙ�������,cH�૊WG� �Ѝ�j�)d��Ϡ�:��[�~�5�lE������5���*u�Ax��G�.ٰ�.i��*���V�LQ3��@q� a��d�<���ԇ#����p�j�a��c��A�0tAVW��-�ı9�Um�b;EЃ��-()�
�.)��ь�*���4C������*g�`
j��?�9��q��(�e�6�I�}T5�T�xY�!���䒿6&�*��Y�4#6XP<������Ol�uL�����/Dr�⥖�y�����e�<8[WVzgaJV���5�����E+���!U��k��	�x�q�j����bg��Wi���E�k����1��_����*��>�of���M�"!�C�_/ �n������fk\d�oy&�F4��dfC�RT��"j��o��ŝͣ�j
v�b_#�ةM8�q�t�g�*�	�EH��B H��5�7�;�9=���so�Ϟ�ڿ�K�b4Zҟ���©m�8�r�����e�)��`�,f�"�n�D&�����x���njg��^�F���ker=T0BT�`��g&�|����O��*�W����4xu��������,
3v�YS����- ���ɥ
����zt�}y'ױM��}���Ċk�۲�}7�D��ΥC�9�.>k=�7o8>ļ2��ւ����)�>��>�ϟJq�%��.9<�����|2-Q������N#چ��Vg�c�K�#�o�ۆϴ���x T-5R������	����D��8��3ÿ:b�h]׏�<[� �f�8�#���୩$
���Ov1M��?B�q�pK��/��6��:w_��4��n<�b��ȑ�����N��92Zoa�8��Ά6��_��m�ܙ}�'�jx��2�Uq�ԐHYS��iI���J��c����PA�RZ�qM����D#읡�$dHW5{.�me��x��Z�uPwj�a�e��eiM�T�=l| �~�[L�.�Nl��w~��	Ie��@��a�<�>
���0E?��tr�W����)y�	��T�W���XDnl}�AV�����f	�*��h�.�gXd���$DO-��
ܣ1vP�3$6=�n�dt���O)t޵��>
���4��|_�o���g==�*�>R{�[�@�h���`�X/]�1�\�T��g��RPi���Ě���;%�,�ع��ߥo~��[ +@�Y>�K\��Rn�1ڌ�6�)�CX�M���+yX�z��G,�4F�K�:�Ű������h�vKʪ�=҆�n��{s6
��J��!_km��?�!eL���Ύ��Uf��N (�m��`G5ԯ�n!��ݳp���l��c���P���B-����׳H����_�񤒦�H���v�&�ca�=}�UǹEX�k�C�e��y�o�Er�Df�4/��8�5�@�(�r��Hh�=���]_x^�*�HZ��ݢ��UiG8���{���p*\��+����rC�.3cãL��:6Ո��Bi��}U{��/�0�������h�j81�{�H��R8%-��� �"��A*���)\$<D�v����_q��]����m�o�$����&���{��ș��z��t��Qb��u��Ļ�!��������Q�	o{���3o���Ӑ��Yl�W���SQE$E��n��>�7�5�--��_��V?G��	<(�z���4�D����/bc*cx��=���:_��d~�rYW�o���g�˒��.D��+���[m��>!sAʼ���]%���D8N|:77Gvx���s�"�	�l������$�	���뀸l�C~�=u�7e��v^ �
-ovϤ�]�E-�7�dD��t���pĮuQ��K� ,9�զ�&%F���,�&&ԁ��kT�}�\H�1>�ff��$���I3�;�P�}�_��-��˙Y4"X�C~i5�JS��Z};��|�uW7���bOx潿�\���-3]��ǧ� �R�hx����ͽ�ЖA�<Ģ]
WH�R��n}�B�x(2r����{퍴<i�yǹ:���5�{�"�;�z_���뭓��!�&Z�V�02JB`Q0tu�=��9̔�U�OG�!��V_Iw�-�x��	��v�R�yͳ�[ST�xٸ�������d����-F���
2�����/���9W�G�����ۙ���R!��P�T�\�4vs�1)�z�.R�����00�����5�GCDb~0F8>����� 
��V�G����$�@�q*.Rx����32Ju�ɳ��+�*� �.J�q#�\A��Rz@_����"R���?>� K�9���W�z�]~]R��H�hC5�B��p;U�c
.�T&�RٵP��3�8�Mّ�}E�o�q���
�k�k+���r��S�,�� ���2��<Τo��zfk��}�=y�Μ4�J �o1yB�_[H�Z�<)�QKpJ],�!^�NϽ����:�Vd�cVY6hǕ��|Y)*�:�Ғ����v�5w��UH�-�ĸİ�~���ܞ�~�]�6���'�CPQ�5�_7m��κ��C�2<m������4:���+�5�?M}qd%�É������6t"x1>X�@mTH�,Y!$?	�N
��y=���=���Br�/9�?l����b��Av��C�����ջ���j~K^�3�'O�|�n��Ggћ����+pCЯ��u$���m�T�c&�#c����j�c�夹\W�Jn+͸�Gkj�&`ld\�K�W�~����
����=������,U/�&�eΘ��w�jn�us�
.��{�JL���S��\���V&%�b�	v�!	�K/�^��x1`�������9Bo��覮��2�m�h�����i�9�
&�E��G�*\��c�`t�?��+�)�
��H[OJ�W�.�N
�R��Vԁ�[�^$��XL�5�5��5�8$�3�0ysS�L�r��Y<y�RT� ��\J�Dc��dRjذ؆�t��Yȼ�L,{��Dx�
��B�~J�h�Φ��wD�Y;��+um7y��p��Fj݃�;l�<N��w��L�����>�w����~4�{b�&g�#Sҏ�H-��ϣ�,��XЊXr=�|��8�� �����A�P�f������{\:E�r���[������ʉ+���0)	nk�{!l޺0�ԇ�LC�N�sC'M�����|1D�:��3k�ny:9R#��ك�����(�|4�Zo7W��çӉ�3���Π6���k|�(��4���F �uQ����n�ΰ�� ���O���a5��]��XO�rZ�b���	�d⢞��v����P��A0X�� _�^�p���ث:2���Z���1�� L�h�P� F�jJ����p��S����Ĺ=����>\�0ZN<�����Ї���*���60����L�6��\?�@~eԢ���F&��h���m/����U�L�g��ҁoQvO\Ze}g<�t	�;�qI�s��J�4\� ���Io��'�t;����sN�n�����:�jm4N\߮�n��
���"2�SzU%�z5{�WaV0�:���,T̩SxX��ˤ��p_S�)��ī I���*�f�~㱧�Zʍb� �=2�H�n�5�@hH8vv~�vD�����PA��L��,�6�Z[���m�Z�Ou���1JＳ;��Њ�J|�Y�����q�qHh��vɴ�^!�oU� �`�l��G+! ٯV�i����'��x�J����չf?�����͋j���u�P?,d��J]7.�6�P�w� �?�~p�E�2Gdn�{��֖�����V:Z�0�Ш��2d0�n�:�y�C@ ,I���]�/7��M�B�.Ңl��Δg�l���K��:ba�����!@&mt�w \S��֣�Q�\�����P�̄�����A�c�ܑ�����Qx����8���T�oά�sHOV�6ީX)_e�Y|1"S{j�W���T>����Q�]f�Bj7�;���U�z&���G��]�G6��ʱ��6���͉�*R���f��U�g��dG����꽮���%����:�P�rc:��G<�  �snڞ�sx���~;r�`���s�肨� m,��\\��ѵ	=���F���o���P��ޒ��U��l�nk��D��u2pi�%���V$�Mo�NDD�|���۹x��\��g��PE���k�yR&��Z�e2����<H.~�'�G�x��� ��ض	��Hk0��Uh0c^Sl��?r4�
�}�eh��H�mE�}-H�~�7ОzAf�i:� =9����7<��Ě ��{�����pI��MCʪ�7�V�b�7��PE@ˌl�n�Ci�ݭ7l3U��:���æ���u2���a��8o�������^^���$�@�M��W)��q<����F7X�,U.���adN&����8
�j?���r|����hrS�L���Mb�Äw���wY�?.a�7��GBoӳ��ؘd�*�{ul��R�e�r���RJ���􀔀&�
3�F���nМz� Lǉ�&�it5�'b���:+�9�tv]����9��1��,N����jY��Sf�����k���� ��H�̮(�9���|-��6b�]�B�M[)lʛ���8{�0/����1����JŐg뤳��#Z�U�\,K�Ix�l�WF�m��">����_�x6���/��я�#��VTƁ�m!�Y
�k�
I�K�d��*����L�ۿ$��L��R���Kɝ������IO&��<��w�5DjL�1TY��"":�.zX�*Hw�E��.�^R�*��|��	�m�_S����Xn�1?+���VMǖ��D��G�w���ؤ����]���İ�����'�����k��o�^Wsa��Y�CΎ�5��hj��SyHM���d$��A �����7v��'ٗ����Y��y��9�b�7��pI2�U��,�V����L�?�$3Ux��Ư�$PD�ȼ�Ӌ�������ۣ��0�G�t��Р����M�љ:8�P�h1�:�����/O�<#���ümDx �[{B��N�rGG�f��z��c�c�
�c�=W�Z 0���$���Xn�w��)��t��S�y
ĭL�m�!}U~�Z&a����A+�wH�lJq���ۊ��x����zϱ֕NzS�N<�묽x�` I��f����'V������cE�d��o:�4�C��Gi�	���U���`�����(�ȴ^�b�M�E:�����z��o¶���aZN��sF�P�"�[�����l��ή-�I���|�*���Uݔs�`���+��/BK���*q��,F��C\�7�Y���Z����pq���Vw�����l��!yd�F)��XN�!J��<�R��O�7����;�+����m2a.b�؜f��D���<`��CLC�����&L�,�,�q�9$�p�A�S����jv[���������}N1i�����{8U��@����q����|�+�0Dܚ�H�ڎ�V������P@�ݕ����N�`��->ؕ�7�X�������U #��R���Twez���ٝ���>F�0�Ԯbq����a+i�C��ȏ�/�E�>M~'�O9� Ӗӆӱ�k��?�x����:Dl7;,�y+�G�C�9oz�f��S��6���Яڙ{9����ˬuaUg�� u:j��0vd������а�F�*�J������?3�c��2S��uɅ%�E�sJ�,����䕎z���Yn)
�j"�
��aW���'��mۄ��V�2
�Q�:h�V��ZW�L*�}o��5Tf���r�P��<8�*��𯙎� �>�偵~E�Ӂט\�8�{&aҖ���є�}Z���؀�╱T���{�Q������;)��E%�x��������3��-5�9K��yq7DX�ĔU5s���W���z��\t�؉H�2������Mt/�s�:��:��������3vJ��x�z18Lo7����6��r.��/��A�Q?P��җ����$C�ڔ�6D[����Q)�g¨��^�(LX��
pו��ө�IZ���&r~���	�x�et/����.�r�E�fv,48Ѫ��Y	��t�.�3Z@�C�^�:��%��e}��!q[����؊!6ѯ�c�"�nt��C���u;�-e q�H|	����Ů��)��RD�ae�!��>��������)�����L/s���=���=I�u0�ހ�t�چ��8ӛ�� 5�op��_m�'�� \�������W�� dQ���7fHY�[�Zc0R��%�/Vr��� Y������H��LrPCJ�´/�dXT3I�y�n̶�>��r� h�@i��4a5A��^~�b�L.�HA�w[4ANY�Z(�A)(����F�Q�$��-������n+Sk���~��������?L^a���zu��K�Y8�Q���R۲WDhQ�^T���t���r}[�P���+�>��&���:򊏶��$�ֿ���\��A8áR�r���
����
��n?]5'~I`�����x�~�W���l�%ޔL���:�Y�Z��u��o��f�ӿ^xr�@�j���3�n��4����*���H��v2���#_ij���Zq�T�3��e���8����'�E]�BtJ΍? ���(�t�O��蕑 �%��mW����+�[v\�d�Y���YȖo,XU+�mEa�9(��*|�4PL�Ï k�Z@�o���k�3���Z��]m�iw�Z�l�H���/6��3�88J)S�."�
FXG�?R�p��%,�[29�"60 ���a��[�{5Nѩ�iz\7s� 
U>6�qđ;�;����T<r~�T?���j�\����3���o��o��HX9�K�S�Sx`F��cΑ�ېdEBz���Nxe�|}������'�QI��VghpJ��ƀ�>�|{�\ס`2��e���m��'��K�?��/���3�������!�䙧�޿^'�5$y�Ҹ`7S�e(��$
�pN{Wd+ܵH(�p?�m~����Q��K"���#-��xn!���D#q�R!e\��=���r�*���xp�O�.�W�I�OD�ׂv�s�Ӵ1ުukSDn�8I���fS�5��,�N�Z��dO�� �F�4��p~�XH��-��s�IjHÍmmu�R+yo2_IM�6Q��ʒ��i����<��q�ȴ	Q��2^F����9H��bK6���B]����m��V b�5c����`���8@e�P~�
��in�`8�6��=���at�-5�n2�"�?=����Y���?���Wġ?ɻ�\���M��#AQ�N��0비�����,��UD�
�(���Jy5Zӗ(.8GM�Fb�ߢd�>��A6\�Om�5C��"��2��t&T���A�	�&z�xj%�8Q�g��0tZ}o�}Z��o�ִ���,g�-Hq���E�V��lx�sV������͛�Ɖ�,+yp*A=�q8c�'�v���5
�۬�����!���E	L��)�"Si��Qq� 7 �b����9ȗ��DF����gD��&����J��PK�P��k�ZɨOV��v!Hy��{E��F�oYH����f�S}+-��38���h�)����ķo]�6��B��=<�j�2<�%��l�V1�(��n�Э�F%�G�)Z{�@�
�,l��B��!?^K.a�}�$��D�o��{�e忦��Hhk��l�EO.�A�9���J�4����tߢ�=�2C��W,؏=�֢�u6�»�BF@���TkEb;UN����GU��17"�� �H��;��I!�zW�4{���,�$�kfE�/y�ek����I���#Xd#�b�X��_]o��Z؁��������K�˜�+�J��ŷTFq�Y*�(�2�>��3�����W	��{�;����gf;�����`'y�I�aY�f��@֫�[� "�*��f�6q��"�"�<%wf��?�	Q,@��3��s��}1�⓲������w _�ܵŦ�_�%|*Vo�qTC��2-�C�7x��/͛V9a���þ��A�~:Iw�Mp�����Ր�:MϾ�7�����������A)��)N����A��9my♍��9g�^`����>�ҍޕ|���x�!�
�靾��]�!��bۆc@�{	�Oa�[�]; w}H��&��|��lՆ[��H嫱ӁZ���:h�;��NK���fg\�^4���06��/��:�d�$"���qBm�{��\�/%��l�F	�ߏ&�3��2��4���f�*PN8q g������bz��ͪ{�����%s�� L0��X.���\��4A��F8��:'Ma�c4����ں�3������L�	
lo��}�00�*�a�;��ʟϹ�''�P\
��m�K�� d�������C�8���k��d�U<h�,�l���v��g�YSL˂ ���0�.��f�$h�fl���3�=m�������Ǒ5eqg���$Y5s%��ذC���i��T&�&��a뉚fΘ{��?A9��f����Iӵ����<%�����澙E�P~b����5�43�0S������Ͼ=%�����Ea� _�Lþ�7�ޫ?�at�U�� ��j�-Ut��ܙp�,��I�#��/�	7ڦ	���X��ݫ��(Qi˧�m��J���32a���zD~��#��03�m���ЪP����*�����M�;A�x�æ�(a��ܙ?.��n8��YY�ÿ�c�P�s�8���y�K4�rF0mj�^�"�v3��	��=��^ȝ�ʦ$yn�n��$���?������� <:�%���}'�f���~��J���v�Oo"��J���}��(K7��й*��j��,�(R�˙��v��葔7��Ny�'n: ,�Z9���Y.y��J+����Ѝ�:�1֯�T\�v�K,KnSK��2���b��#����Wø�#���2^���bF��rl`��Lo��0 �f���ի0侢�-3�B����N^���UQK�dS��8/Cr�q��?ږ�q��BCǤ�C�+읕�cŋ(��HD�B��"Q0�+��������1I���-��^ i��PBG$/�E��dٴ�����FG�(�F4�v�8Μ.�W�"4�a���)&�A�8�9�O[�$&��0;V�`��ԎW��v�q�<���8��Vפ֗fBȋq���H�P(�����.���}\^r��X!ݞZ�n3�8���9ϐ�44PSWZ���@\�Vu��w&%�T������n|1�*��*_-�ܾ^�P�]a����2�')ps@5��x  �6�����k5o�"R���?G,SXd{�E�JO"�8���m���|�?�6��>��=��jDرp�ב'�M��j�r�d��ͧ�����|�}�u�q+���|�)d���Dqٓf1s�m+[�*����SC�U��Z��0?���ǫn��}���Co�p���K��������J�A�B��x��vofӂ܉ØT	r�kϑ�d��ԧ��F�{�~���i�S�$7:�<G>���B��ߠ肦���Kp��,���l���>�] 7e:��L�3"8G�6�BT��w�x�O�%��g���&�g�X�{��f��F��3�0�?O}:��ʉ3ٕH#w��Ɠꧧ)���l����\p�_h`�	Сf#<K �`dKm��c���V�k^X�,��BƂ�O_��^:�v��j*�OP�/��zg
�C7Q#=	r�����qt|I�7��x��̵a�eO�VOY�z��_`R�o�	R���z
� ���r��t��T��+$0f���[��R�O���{��0��AjGAc4�!��7���t�4/k�N��0g.�R��祈GC/����㥸�Øm��y�i�v������.�MG��d�_o�mDkE�ZAGH��&=
�ܮ���>x��Ŵܨ�o8�1@�̸�G�i7�;�T���A,{�al
����O��$'���ә;�dSP��k��,��L�ikr�~�i��1~< ��6�eP����v��75}�H�l�9��i�Wzr=.�0��oe�)��H���&K���vxy�����a�������]�����x�ҭ7UH� Bwm�d�$��u�h�kA�@�5�(�$n�-���j�A��6�����qO����ذ�-�-���n���5��g7@�C�֎��iy�΃���C���0�>��^XuQ,���ы�Oi�m�r�7o�� ��;����g��j-��8J�a���n7F�Z��7s��:\��k���G='Ձ�~�������ZB3��8E���мcډ�e���NŮ}34kOv����&y����O��b��%���&�.@��|'J��T��Y}X�A<�E,�ye1�#����#��3�:�x�F�B�|ܪ+)����,0ڼ�6��JL{��eQ�;@\r��zg�}ȿ1�E��""��O/�o���7�+r'�&ͻ��"�����M/2���{�>(.�n��=��]RX5LV�+s�a�]IZ�P,Ԇ܇Tn��\�a�Ҳ��N,�$���>^n�$�Q�O�$K���]`!��:��U�W�`�!¶�<�n��Em)Y�i��g��Ep��Q���x/-:�m��u�)�+�'���D	z&��U�E��9;�!��F�Sџ�dfN�L��?�B#�>l����39��1q�����,6�sj|EV]6ڄ�&͈ck2�"!�H���x������	t�;����eΓcV0N�V:j�HJv�n�`��؊-m�b��C&�s�Ç ɑ��:��vf,4fp�ݓ��]8�����1��V��T�����.dӈ�X�@��<Y`��#�,��'�u�s?�z1e��8���L��IQ@�����/��e	�v�+w͇�u�{;���˵+-t��v<�8��n;D�E\����ZQs;�S�N^xa*f��B�~;�ŗl�)�>A\�~̰���ԭ�rך�'[�Z�tV�bz$���y�KZe� ��+���"H��<�$�{nf�$��T��Fq��P��2k�z�q-��]���`���N�)���r�ِ9��|U���`��,�'�G_ZW����)��q�;�6%����N����d^�������g�0
��K��=��[Fϖ����t��n��q�h	�h-Anf�����S�ŀ���뢸��]�uin� ����9��^52�9��'~��L6`a���F�!��p�!�� ���n!s2�.um��B�V�|Tu�$��6t?�s\��&�x	��Z'�L�	���Ȼ��J)�=bc2�g��	��i�����Q ���-�%A�3t�O��+�1�O�4���_`Z2��S�o#����>�Α�ǆ��<LC�Jvt
�	1o�����#8y/	}�5��e�L,�mt��\�LঌN>�:�_��A���8�f��������z���xdV�V�Y��޴5Z��65_�y\E���+�t�Aa�fh��؍s���u<>߭V���3�j��蜡XN�$�%��^�F<P�C%�a8��W^���'��]H9n.�٧䚐d��Ňpy_��X�6g�gѳg���qZ_T�{_��;���1xV��o"!��kU:���A��B��(W,	�<�r��Z$��l���e��Z�*���>���"h�A.�$�Ӥo���g����Z!�>Q�ov|��/�Sb.M���������,�2ِ\�n���]'^6�#�B}��m+�s�{����$m:ӓX��6�(�<�
�3�Y�$g�P%��O�i{�S���Wp���������w�$������4X]��!��Z!��U,E�g��n��X:��6�?W�g�b���y&K�5E�8*���q=Ytヘ��B�uLK�[��$q:8�o�k!��D�L�;^�n(j�3�n�%�Wy��w u��+�Ń���L����4gIS�����(Cu�n(AsX�}�O�8Pq3	�!R�{���CW%n(T�x����P�㓡��o-[����T';�0g��Y��� � �f�*��B�U�9��#vg �W��?�|M�6s��7C��C4�R<n!�"|�I�J���dI��E8L�+$�Cٸ���|����(���T�������$����D��v1��3L	���bӗ`��}{�I�YCr�G�Z��_f�����9w�/�+P͆�X � f�A����^��fOR7"បV*�8@	�W�O	��|�͆���=а�^�Ƴ�K�u������6�'��w��_Z�0�mu����#�XD�����t�G0�^����d�W�Y�!o��f�����Zy8��eU���q`���+  OT�7Ȍ3���~��8F���8�y�`"��e�,|H�s4eZ�p��a��@��HNK�"���)���?���Dk��O��H��%�-�Р��˵���i����x�+���&jq��	D���H�-h��� PM�>��� c�{�5�T�]K'~�]�r�o`M�\��� ;�oh%N�ܱuU
��T%(dPCxQ9ܣ#����Կ|k��q���^�[O���zoRU��� ���w��8i�`����2J2��VťV�N�I�bB�z�f�B��e�Ջ��_h�Or��Xg��5u_Wwo�P�<k��*����-\5�]XQ�L"��h�
A=�Kny�37i����kb��TL�^���J��
h����S�:ј�dd1fK>z�j#���V�(b����yr���
��n���0 2���bp�Yb�4�q�Bϯ���,�O �ӏ�
Y;یJN�i�&J�ҝH����&%���Է��7�2��5g�;�6M�-��N+��ts�
@GI�����]^@Ka4¾��s����I��	G��0a�h*��v�����-����C��<�x��M��qP]���o_O8e�ĂX�aБ��E+����x�������8�nVN��l��j¾y}+��9���;h�o�&�WR�YM(:��j���X���Q�pM.7�Fa�Y/�n$n�l ��*Id��K���0�.�F��Fu76�:�f���C��,�N3C�[ÿ�q��OP�i3���#�V9��h,�\�ݜYuo�ذ�zLЏ�d���R'�H���Q��0U��A'f�]M������~���1��֣��z���Rn�L�l����u���\��~�5^ʵ�f�'j ��x�APA���,���R���O{O.S���4QV�@3&0hQ��P��K�H���W4$8\E3����r�g��Gm=�����4�T
H�mEA�B�URWk�c�.�,LP��9���D��L�2��4�����*�"�s����p5�p�h��?����j���"y/����|B�fN�}6a��j�G����Y�R$R7�uF�q�׮�X���npPp+\��L ��G�M�d��	��N1K��z�a���	9s0�k�8� G��ԃα��D���G �!�X%m&�[h������T��a�w�&�0��T׆�"P#�/�h��¾`=ZS�T �N6��_%��A��7?S1�uJC�����w.�7F|�q�[}��d����(�E���Ms9�I���`�{m��$����2'o-�H�D�δ���GkP5�W��s87b=z��Y�o���=:W�Eg\[O���N롞,�i/��K����v��ϖ�~��L5� _JX	e|�O�ݾ����;���W��ˊ���J��}�/q@z�6=�2\��mYU<�uV5���]ѩpO���8A���~Q���ڿ���d+a)��1�oZ�u��������{��<�u���~����}B��'`Z?��	�B���5�-�7bW�/Bl��K�{�y�	wAk��n��k��#�UA���[bͧ���F�F����tU_gЗϊz��G����@[�>����^U;ܲ�qR�H@�XJ4p\s<���d��F��2��<j0S�H�����p��-I�⊬=bMS�̂(	�Z�Ǥ��Ԑ�d	{`�Q��4Eyc�o��q6{%
��������ښJ+�Q#i���l�C���ú���7�[�i��0��"a������R�CS34{2�|h��ݬL��Ь(���j]w
�J������d��;+B��ƚN�.�N^�x`�=1�!
Ȯ��ftZ���ސ1b����!^*D�o��2�N�o[?dp� ���T3f5�>qz]o=n�V�L3��}�n�f0�H�ц��Cw?�C(Q�6]z����".�v�WGʜ�d�"��o��r�mYPA����~����&˒76������$!�~����)Qї�&�u���Q�V��L�3��R6ȸ��Z%We�0�溁��7�W[�?�t����57�!ҹ��T�U�N��T�.��k�27\�х�+F������Q�Sy^�p2it���8 �zeo����=��J�V;|����~�
τVj}��=�Bw�4S�q���QQO��>䇪�!g���'���K�K����o�WY�����*I�Ҷwq۶W4��rJZ��.��>=��v��#N	Q	�MV���-M*�+[,$��1B@�>{8���6�i+��#�32�Ag�/��̵`�_��+՞NS���6�"V����f��ޠ�ط9�a��S�/"X����*�W��۟�S+�|9��%��vO�첒gUm�ػ׈-h/Td��O���1�~0gP����i�QG��fElݖ(��'$������9���1�m@�J�ᖻ`��yn�oPM�����vSw�H礍N���@8P��3�-�Wy�R��RǊ�h,^Mgu�ȏW��e|ݵ܇!q1 �=Oܞ�I�Á�a ��kD&H�g��hj��m!�}�h�_I�y��hE��9��-�^��g����rN�r��r���A���j�
�r4�<ڷgK4�i���&n��)����b�җ�I����Ef����9��r�g�oAD�ʛ� (.��_2mN8
�W.����qۡ�BA���E�P�9: �I7���j;�`���;0`\Iyە����6l@��_��a�[�h̻+�����t�"J���Zgj��ց����s�8hB؎�c��?��]x�GK�u���
 ۭ���`~��{4�B����/@��S������4�s��7�'�n��nM���j�)���U �\���I�H�T��u�3I����G ��Q��������oF�Nض{�.��`�b���c'��+������1V� ��?�4�P�h�Ւ���v���G���>���/ �D��xb=�bdB�L�������Ħ1�̐ǧa�a^�X�v}��<ffw���d��zJ�~�Cſ
�Sҷ�0�L ��#�d�*pyO��76���#�Z�)�)�ɘ���V5m�w��Gt�KZ�9kg���/N3õL�8 X��Q�g��N�z��x��S�a9Z��`o�M<����t���-�劑U���;<A�:$^��l_�)�N�1�,��'ym�LN#I0&fM�3cW�mar�4m\����Z
9�Δ�6t���M�ư�&�� �	Z������i���S�?(]�z	�h��ʉ�b�ז9�><�;(>��W]��xY<�xzU}���1^���rS��c8&�����<����l���8܂8^��_2�3�~AE0��>��K*$� ]�	�VZ��ao�/F�����"�Q�5Ã.=���N���ϝ�|�_�MZ����H�F2B~�����FӼ,X���@ZW����q�l�Q���WO>�|����c�î��dj��G��?�̜ю���xq*_���n��xx�$�Ҕ&*��x�RCrk�\�B-t���([�/����q�R�,�����Bl��X�)�G�K ��Ҫ����<�Jpj�2kE��TյC����ϑpS�Y��Qt���%`�`��NHf[B9&��z��xͬj+�Oc�3�D�4u����?�����t�EAH�������N�������"[w�g]��	s1]v�X��zs/�����1g`�N�܇�KK��;�7�EO�h��.&s���'8X*2��{��D�&o��*i���W�"����s���F� L��u�u�������ХO$
)��5� ��#��[���Q����c�|����0<;��t��UG��L������y��앻�eY!Ne�� �U80�ɍo�?���F$�I}��
;Zs���k���7/�4X󸝍�WҀ\��`G�+"�m�H����S1!�j"u�����B�@9`:������V�89�����Al)��w��Z�����Am�ɺ5��ꍖCG���r�����C~�Ε�����Q@�����]�\K��V9�w�%�^�op�Y�_��#J��L�!�}�c�6�E���W ��L+���jU�*���f������u��5&m!�r
�"b�D}�ɸ�����bŷ;��6Z�����'�y�Cq���$��zY�ت�b�JLFmdC��EB=���׎�Ӕ'h��%�T�A`ZY�P���Y��م���6�Қ6�� �^��4�J�1�������۲�o�d��8ع� b��4J�r*��P�)�{�ם]���^5A�<ĎsU��ɬC�W�`��1���I�>`v`(Kv�"^}������x�(+E����-mN#j1�E��뚹���������n�I�ٳ���pr����>mqq��x�2�ر�9q��Ь,'�qt�>.b1�Ҡ�1p��|�;1
���|�ON���R��v�],'�yr%���oU��!ː�tA���LT�����5}t�����xBq���ik��wQ�H��(I��I��s(�)�t�̌q!�������)Dr7Y7���XS1l���~�fH������y6[\=`s�7�I�
%�P)O��B����	��).�������0���p�C��W�v�J���Bj9/� ����S�ʩ�ڞxK�9l���u��w��J�c_�����&�!��������#p�R)�^�f^f>�e'y %M��`�j�2�i�;���U��+a�����-��S��0%\�<n���r.��ib��J�&�J��.ו�bpJN����8��CFL`�zw�&�e*��^�d�wz�6��-�W�	��nl�2�;X���p��@�ϋ3����Q�T�F����2��H?���Q����8Sơۢb���E��9��	T�'�`
�I�n&�̣��JESL���7�=�Ќ�^j�#�  ���w]a��ꍒB.wBix�8�Pl�x��	��b�bR*%_�62���'�#
\� ����s��?t�WI��|�	7HC���-=]М4�t%�6<�a[�M�;~��`�_���Z������<��SHԏ�OQE�4R�i�	��ޟ� ����y	=qq\m�C%Ǧ���si"3��-L:���)�s� �b�r	m#�C{@��F|�2be2��/Ŝ���b.��q@�(ҽ�S�{�A���V����1��sWQ7�-��F�4w�&�0\�/�o�^���L���;������h����E��Ϩ|<�aK(W,W<��E���!�f�v��~����`���c�Wxw�Xf/_PF����O2������+��)��}~��9�h8I�]�6����e�o���x"`��� a�������B���Q�\x��<����B,�m����E&5����*�z1�I��(�]Fz��(0d%T~~���rƣ�$�ښ��l�q������/q�0�KJ8�
�=�ZdE�v�tw�ra� ���q���g�*^���Cږ��Nm����ז|�2fz������s1�8[ ��5�;�})��04?�(���i���kAD�q.+۵�H�pͨX+;P-;\��g%%���d$6'�v~�+�t����+���	����Bqvw)��'ō��ޥ:4�$ 8�흊ÞP�ϊ��bn�_wwu��wt�guP�7w�f��]i�>u��q �]p�tUM�Pr�}�gn4 �c*����`�YK����.
Vnu��խO[Zyd\�����%��J?��X��� �ނ��
a���_�Q�&r�n��ݞZ�JA?a>�kHů��"w����k�U	T��k(2�Q�Sʅ|:?��W�2��4����\��MZ��N� ���Ka��2��+�r���q>P�:���CR��7�,Nk%22_�Ok]ov[�3�!K�	<��|��x��&�!v��Or��P&�R�*p�~Wx�Q��NI�V����ܴ��t�o��y+Ccmav(�1o@Q�8ur���o0���Ҟ�0��d~�BƜ��ߓ���W!�-�?������g	�r;��C��E�/���z�~:E��� 	�vo�΁f3K3C�����"���޳����>��;D5�>�����%�!����4xo��^���E�����x�u=�07�i��5I,�6�c����UaW�:���/��@����~����n������FI��e�hhFC�H�Vk�f�lV�+ZX%nn(��{�9"���8��WY�v'?-z�^u1�KqZiͷp�Y�V<�ޝ�8�����2��U�����HT1�AlQ�;+����։Zg��4�|  ��������J��������)���W��ά��q�6:��v����2M�o��v�k�t�,0d�ԓL����<EW����Jn� `Sl�f�Y^(���¿y�z����f�j9nTnO]]������c�\<�x�#	Q��]�A����(B،�yT���
�����d�*�e��b�?���)���α��jDE(��|�agm�ڼ�����a�\#�k�w�n"ׇ�G5�� �Va�t�4�O�/�N�ꑒ Z�q<��]˳��|/j�Tu4�qe�觻����Ԣ�D����:�ˏ�ɓ� wf����O�h�C�EW�Ӭ��מ��8�����?��5#s(B�i�j��4��VJT�#9���\es���SQ��YP�����D��<�NDbZ�z,�4��pRoFV>�֠q�d��>�/I���]@�v��)�D����$�����LΏ��g	����!@a�Ak3',���b��eT�B:������}2�=�*e�#\Q��}�lx�����"���7~4RUa��dm/Vn�L�Fl��Q��_r�%��d�cj9g��Zߒ+@���|���{����kJq"r�h�Ivփ�O���D�)��Ƨ�������o����8�6r���w݈�%)k�	y/�:%|���z�?)Q\bC=d�2�~n�o�;&4	���Y����$�]�HɔU��~M����̃3v*����J�=�����1����L���҆��PX�$q	d�����A�f,��/uN	S[�e�)�)��!�m̟8�t����bsdW����� �]HV��힗j2#����l'��,��P���|�i�)=W�s�д��`�Wņ�i�iϧWAk�i�x��ym6��2�SdJ�h�����tQ�c��q-5f���ך�B�N�#��^Y�)�x4uE��U���K�W)���8�e,���?0���L���I��)p`r��X�o��100���?R�Ԍ�?
��]M2Y�ڛ"�.�x��-�<��u,]L�=�`��)�����ˡ:u_5���1�%p���q6܉���"	�&&��N�D>��nxm���j�&�Ao� �G�'	�3���@���'�c��1�3P#I3�@��7v.�}��g�i8J(u~��i����)$y��x$FM��i��Y����gS���� �=���T��%w����!��91,��ТR�{�ArxW��m1?�х��ej�=ŵ0��i>N���-A`!���}{YM����@9�H��N;8$��,7Ӄ���F!�VРKJAò� r)��V��FVj���D��S{��C���+��{1�""oÞ���x]Z�,�Q��,�h�&��$��ɵ0*7u�o�ZՈ=;'��������㤸$7��p["Y|_��p������gNf���)d��+����y9�$�v}�ӷgg�w��7��C������}+��e�uU��ϗ��yX�;�#�VdֺK��GF��"j��4��էC��o���̌~h}���B��}��|R��¬�R�Ἷ^s��EC����ؒ$us��3����ȻX)!�h�0��Yiշ��]�u�^��	�����X�t�B�AнQ?�������BC�C'��gRO���}guv�Dm1�Nꘇd4n���i ^�L��ʦ��98ۜ��.�XD�\��$�'�FJ�����.%k����+��hTO@��,�����0�V�8{heL���6�q[G|ؔt�y��>��W*/EmF�q��Y�� �mI`��{�Gƫ���a�5�oֱ���'�޲�:�����Y��E5�	j��+S�����
Ǿ����ܩew�Ջ�>k��r�� �)��#2x�D� =�38)NV��>M�0p�$�S�ѝ=�~=���=�]��{	)���ҿ���c�	Fp����C���& fHt���C �!�2h���o�@����b����{c���z�	#7�t�,y�!��<�)G�����x�=OrΥ��A�tj�4�)�<�%Ə�����%���վ�jm���� >�{�
�����P�� ����,�Cx��J�S��5��mE�LN��8_��\�E��ЖĒ#��2A��%�ot�������2�!�%�Sda'A��h�o�L���~f�=���+�	���� ��l��*�:V\E]ً�ECV�u[C��d�Dy��1J���C�.^?R(9�87/�P?�CFx�\�Q�=^������9j�!�d��b���O�Ҝ�F��t-:�g���m��V0:u�@��ʕ���Z��j���WL��E�C�©��˾�!��M7��D�(�罌�`�a�%�Ҵ��e�E�Y�=�PE]ɵnQʴ�����Q/���=�$�U���
�c	˪P)�z�`]x���6�A��9�eJ~{�x���:�L��_�l^h�I��\�LNȘ��K���T��ؗ��QS9�`~�4������,���-���Z\_�琅cǨ��^w)�"��N�k��W��,����nf�	��*?(�|�}K/(��E�����P(���	�+X)AC�jhEץ��b����Kӟ�v|p�"%�@iy��WK���h��ۣɘY�ۆ@:}�Puݤ�c0�<���j�xI��#�X�k�;F����|�����r�.yWT�S��6�23v ��r�Q4�R���G���Nb5�|%̎�6�_zQn�T��$�fIP#:�8T��� �e#1ɱ�J��"�c����'ibZtT_;}��c)œ��͖���ϛ�epP���s�'�%�M�ޟ���KPt�w!�'w).ҿ��e�=�|Vfm����A��=���������'f|�z�x�����o)��7� ��?�k7z���լػ+�w�Yv�:C��]�P3�g��x=L�w$�2��2޹%�:�������&-�"�W�aB-�@�YD�6�^�I��[�ly�@x�Y^pߦH�Z�
	��O��A�����F
]�Qj_��B���p��[��jj5}�w)��&9���ޕ5�ԥ��'�Zko�����n����(�om� 0ko��Rn�&��A��}ij���`��G�U�#&���RO�Q�8��ȭa^f���-�Z�n���:!q��,90��'q1a�e�Ŀ/]Z�I��f��9�3B0���+(��������X�_e���f5U�ߟ.�
^>�%r���[?4�_��"�GuR��Q�� ��C�0c��{�%�o�wbw�1��?�T>����U�ڪ3 �0�^Yh�m���͐�JF�7���0e��(`=�!|�o>�����Ȁ��kr����ϰht�U�[-�#Q��^���t��2�����l\�~��z�(fI��ɪd\1뽤��1ׇE�,zD���ӎ��W�f��v�'�:��鲆�������'��Uu������X��I�[�թ����C�{_�<�K��:4��T���֑)P
<�o#s��!n��'�yZ�ƽ��p���A��w��3�Bv˟���:�t�q����U2��\�zTp	$���s~ZF��40)E�{O:�郞D�8m��\^��9qͤ-� #��p�/�ӾYH�6�Os��V�[�@8Iս�0zEH�nÈ^xہ���0�`��ɞ_�ji��7l&���2�~�8;]���d�Ƃk ^K�����b���dn��6$f �`��J�Nk!��bd=#��<m�H��D lI^E*f�;^C�+�U��u�����R�_���~�<��!���?�-1b�����[P�k���y`[�0��@����q`7pe�#I7$AWTaؐ_d5��vҥ �=���i2P	�"�����T�2��"�[T�9S�UU�'O�J�r<�&]�Ɣ�p:b���ed�����N��jz��Э��l+�^ޣS��ڽ��hʱ���L�$�
��m+w֍[�*��%[���R��r�"U���+Ut�M%؛��K(����Y'��gVP^���vf�4�휯��{���e���{6����m#�C�׫hq0�ɷv�7 	����gs�e�sI�鴟�ౢ	�C
�t^�J+��p�b�@�B4�$o=8�����4=فhp~���XSgS�B����7��t��~���Z!� �AQ�z�Y��K�A���m9 ��6�H���� �f�ѣw�2��`hT�Wd��Q)����.k�s��uN0;{�[-���r˸d�4��V�����;o8U)��r31r>?(�zI�Zħ}db�
�``����ʽ�64k�?��O�2�)�΢B�����	$ �J��	NOQ�
�z\��C!i�k�GopJ�P��3Y�X��#����!a%�T;o�f����fI�/bˈ�[��ie�n����E ,Ix�16	զ�J�^��tM�yC%z���c�n�H���D����@Kc'K��Ό���W2 �l��ŀ�U�d,5v�\�N&��~K�R�m���)5t��F͵�����)��h/�f�0���]��/�*�=ɏ����{�C��.����Y-q����¬�4��8t֮#&�Q��F�Q#A�d��w�i4É�>5�2���a�[^`Y��c9a��۞�*!�����)iv/��&��XU����<0b�)ð�WL��h|fyDj!�L[�8�i���+D׾�K����u�<�Q�T�Q��'���B��h�9��`���n[H���ܲV����#�5�q�[_P�Qa�6)�T�6l���ի��P���
+�g
� _�����VE�id6;b��ޛG�� g;2R'!�L�P��F�"��K�|����D���&ބO�������ȾqUPB�Fpn0�F힦��sOxH�.cr�x���:���B"nؖ�l���IM �m�����k�߫��=���ҍ�aԈ:�Z�#1�kP�v�C��_n�q�r�|4���ƿK���ǽȚ[�l��N�ֽV9��B1�},�{/�	qC�r���gZ��f��:tP�*�����Z�ż��UIs��+�ۊOǼ]��¥��7�.\�<��&�Rr)j�@w�h��=fFl�N	���4`��j��Eթ�Fd=�8��k OJ�	y�.�l.`E6̉K����e���kQ��@1It�_��h��Lx�ƈ윒l1��l"���}Qk8���rQ¶9��b�Hc�=ҋ��)��uϞ�~��=��}2I��l��I�0��t� yBg/ݓ�|��N�"7Fe���E]z&��ys�n#߁�[�HӅ<�]'ٛ�4#n�F�z���ڗ��� �I��g�[T����br&[��}�K#�MR�͆��PM�`m�+E�ᠽ���̵$����?�WS[��4��%��֮(wl�W��g
������{�l����j
��Ҭ ��9r�O�%���V��m[�hɈ��������	C��YÊf H=)�>�ޯr�X���W>v��0�?�{(�EI���}��i��&#&D<��������l�1P�P�_KAn��3�L��z��{ѳ�\�jO"��X�:�b�u�o��ZuŬ������4���8F�-�\A��O_)�,u��lA=�Ƌ�;�7��,�jY�z/ �*�o��M�bL���݇]
������c�,����r"�\��~EɚU7�&�uS��5����ZvѦML���e�b|�:�ϸ����q��UN*����6�ɪ���/�?sk/[���v�]G��).�w�/X~�ܩ�l�| 8�㷱�3ʿ5�[�״]��n��;j9��0�I��O�� �<������;.(�	:&6��,�~�]�f�r�7���Np@Wu�%�T1�aKp�K�z��Q�ǤH���*���$�]�L'TAu�^뚢̳����Ej�>7��IZ2�������m �F��%�S��$\�J)�dk���zE�WR�"qh,���.�+��mƅ����w_XB���^�&g{/����F��$�'�\9�.�,#WI/�����Gћn��է2d�H�TPh� �!�q�d��=���+������9�נ�ޓ��	�=��P�~
d)i	�Pzh���̈i�Y��G�����`h3;.����O�cY'6B��K��a����T�%LSΆi�=��i&�������K��\�s���'{˒3 ]W�\\����h�:)����8����>�/Z@n��������5�����.)"�"n�Q��+�����i-����2��O�Ț#N�պ��w}�<��}U��
��^@�Y*@%�T�@�w�.��j�6LY1�q�&���Z6��rGun��uG�����;p��[R���pz�5����>��T�J����A`��*�z��"(�P��ړ#!�"�5`J���čx������Y�3����8D,��9]V�Y:�6.�0Rb����{ҎƱ�+�6�͜�
8	G9#Ufm���3w
�-�b0��m�E%t�ؔ��M
�� ����`żl�z ��t��=e��Jezr�B^*Qښ��&ǹn�O_r�H5߹j�g{5x�\6��g�����#|�%v9���ǊDf��a�qf��L��F`��n��7��W"T�� Y{�sKj^f.�JF�!_f����ݑ|�Z/��M�M"6���7˿@�3�7w{�!��.�>\�lg3��!��ՉX�Ȋr� �����(�X��-h��3a��Tc)�Y����T���z�b��.#3ht�]SzC�pe�}f���`F�g'�M�|�Pt�B�*-a�"ƈo~i�B�g���*R��o좷��f>�o�KHД�=|EGQ�oۍmt�O���(���:"�P`.j:Eo���_^#�t����ߧ�G��HǦ��1�j�3~M��I#�*Ql�QGGZjZx�4��>�!��c%c.���(�h#�+�oI��XɁ��W�N���r6����XV��񒧤gz�mD��f=H��*�j[O�|����r@�&#�����xđc�@-15���Pm3KZ����9�\�:)6��7��E|_'
s���(�k .M7e\�ājQ�h�l �4���k7�mf�)#;g'����,�ѭ��m2�y������i����+�~�w]��mS�ۮ�^\��X�`Dg<?V
(�n*�>�s��!z�V4V6�à)p�@���׬rtD�߻1!Oן71�vCRF�c��:�#  n�s�m�|j����D]�J�C�u%�U��|R�a� �Ķ�ɱ�;���������JR�m�@tT�w�rL}M�Zbr����3�2l!�v�zr��$P���oe"r��˿�2��H�޼�,��{7�[���3a80�Ph��&[4�����y����� �C�X�M"�^u�7Y��)C�^��9mh2I��ŋy.dV���j�s$�Lg^>�f�0���7t���S��z��P�s�����RTB�1G����'d��.�3M�	��U��)�9oװ�0~ɓ!�dCs[�^;�����$#(�ٺC� ]�՛9ţ6�G��a�)��49��2�;��%�5�Nw�؇R�[���p�2x�]}UW�R��b,i�b����i_I��RV�s�/`�OJjzOm��IЍ56���hI�6��7��p�\x��.�>�j���$�#�ܩ:+�'��gaS�K[G� �,nm��&4sD������)ۧic&�,���(H�����8�l�u�Z�����!��z{�	����ݐ��s�s���U�r����z[>7"�G��w�&)����3A�~� ��$0<��ذ�)t(I�G7pN$>מ������G�����إP�a�{Wp��U��a��u%�-E{�L��@�f�e!��7�@PD�"m�����@I�^�D D�b�py�K-�K��T�����c1�fw�#V֡����	k�h[9�#����d�)�7�i��%0�H��b�U\�G���5�����2��N{��mL3C��]C����=6���?����J	_�/����7ڱ���rG��݄�'I.}�ٖ�ܒ���>O�T��(5�m��Qqo����dS��,E3�s�H\#���m�a��q��:�i�U��C�Z�R(5y�a-gY>��ŉ��8�d��3��pA�E���ܭ�XY�ܩs�����Á��'�vBe�=��|7R�~�&(����I�RrP*|'Q��Ui@D߽q�����^�
g^�6�,%��Pm�ɞo�-��Sx� �=��	d<2�󙟻[��g�gr2]��n��w��ُ�'��"+dnl����}���)7)�5S\<a�!V�Gs�O~�Z_c>����EP�W�B)���|�u)ݑDDR�u�Likꂫ2���vujn9�9�k����Y ��C���DX�XH�� 
2�1rdT��#p�MѦ�_�M���&��8;Wx*���8��F��ihR,�{(L,:f�m�q�4�gtz��ܦG���!KP����5��?\;C��:ԓ$�3�|y�,@�j<̔}�X��r�qޅX�w�	I�uf������^������5Vi9�/��g�ِK�im���L���}Hy��}x������c��qA�Rr�B6�o��[�W)�g����QtU�)ʶ�|(pJ O�����ֻ�X��^��Q�;bw=��r2A5y�N��	+�%�|�C��ʾ!��׫�e�_3H6�>$+�ZU�"" �l�t�ޯ3-nw
�dI�}�y"%©`Yu�l�q�p�:��k���v�=և8x��?�p�А��������F�Y7����p�2�)�?�M��2~F����=,y�G���ɖ��#���������|+(��-�!�Um����T(?��`�z�j�-�;�=�J/ʼx���;Nm�>�"�Ӑ؇.\�K�+���h�*�I���1��Β�0/��}Dsyn��%��p"����Ӛ��q�$�4�SxY1�l1(��r����������T:L��P���Z���M��]�1	�N����,�y�P�P�p�e�a��0v��
bڵ�����oc�撁u:�/�����}z�L_���T�A��z8�.���$G���i�-*UWcY��0yV���g�Ϣt��Z�3<�<�{fzG�f����n�-fF���r�.�0>�f�$����9��'%z��6k��	���|�.�bA���Y�	�!Nh�1��d^a��!~=�qοw�����b��{���,������͍�	\e����J��,)0��3��l���U-�
�����<#�G�5��Õb9Q�[A2�X,'�ܤ���m}S|�H�?i����[ ��x0o
gA��{K��)�Ww�dB�~i����~29��,F�pNDe%;\�ϑ�U4��^$��O�M�P�8��3�=%�+��b�n!L��v�  ��&���[��
Yn�Q�.�NL�a��!E����3�~|�Ǻ*���:��=&���S��ޕ�9�}�KZ�0�8�cE�@r|&M�m�UX��J�W�D�ƪŻ{l>Կ>1�4;��.ɱ�1�l�}��_I��v�Dq2�ums���ֳ2gyZ�"��r��Q̇�JO)���5!��Zy�TAR�o=y�ګgB��s���QfBî�7I��sz���K��ӻ#����x*ovD�7�	��PW�eK	5�n��};��U�qm >���1��ET�7^Ǹ3����C\�$�c�'FQ[��'2$����B3_GtbUC��L�ߜ�r	���-�ÚI���*!�t�Zp<eJSU�(�K����8cCg����b�yK��_���u�$āh\}�u��o`.�o7&�L�n%=������/�?��7�Ò�E��+�
���|���F�~t��5x3(����bTǝ�Zt�b����^�C`X�[Vb��-h�8V�Hz�M����ݱ7(��)��vc���k;F� ��ׁ���A�5I	��KTB�tP��I_��B��|�+AK�xAQ
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���nNj��%�A��W�s�3�T^�/���%���Iw�|4�G�Sˋ�Ĥ���r��o�����*�����Ի�0>�����v��� �v��Vp������^{۪x���0`�+�R����\'�wo٬�9i���d7���{V�������fz��0�=�nۤ3=�U��l2�4��0s�g���Sr���2�(.�a�.�ةo��#�3�Y{��NĢ�GgtX������5�Ht�9*��^�TLO�B��|<O�����0�,�硈�S"�ͯ߸������u4y��4�c������4v�_m�fX�T���fޅ��f�V1��>��-\���3�0i� �Z�Ԕ�Bb4��?9.>^��,��y�,$��N'�>�j[��dVYV�Z��qj���  ����#ãz�F��?[&8R���X�/��(nL����L�&��������pW@��Ҋ�ހ�|v��EU��[c��)w��`���(�Xޥ/J8)�E��9$��Y��2�Li���" �2H��̩e@�l��8T9�q��/�\���ioD���"�����F����*��RC����޾�O4�o,�&�1\�RK����$]jh��e+�S��nFT�$�Q���%�EOʯw���O(����<�����|�Mɡ<��
�xL�N�M�~Ydm
J�'�� �?CC�Q����h�d���{^%����t��lc�d3�t���>�=Y�a`\b^
����,Q=�S�GG�b� ;��r(#��9cC��?�T¾(�eGfFy,	�:�l���M�cb��}90<F]O\=K^�*Y�AW� �%�.%j��鄖S��/��.������ą�Iw͓񅃨���2��ڴ�8y�$��'�ZObK�`�o�d%q���\�vBc)��c�� � E˼�Q�(!ܭ�}l��h�F߆Stg��oĢ2�$^��]��F�f3+;�S��0L��4!|M�ND�0��7��4ޟ	1����>Pu��T�h<le��o�k0�4�$�J!%�ծ�(�0�r�A����fZp��1��n~? U�ұ�W�>�򖃽�p��K���N��n�ȾQĢ�(Bm8>N�S7�h�6���upF�u航axcpJ�7ܹ]%����0Iy��i�z�j��O�j|��xd��>��5��߾��I��� �&H)���BKLH��+p��+��[W���2��=:��ƃ}���������Jպ-�ᆗ��F�y��K�\��T�s_�gk�,"�������2�q>�F �E�)��R���;�un��J���/L��ڴ�Ř��XU���tz��OӚ�2yz�����M5�zM���y�^�|V�@�t�4��-�6�r3@�-k �oI�_��zk��0+00
Q���;�@M���`����N���6�d�E��2e�4�� \sZ9ƞvX�3BP�ǥ���t�{�|ـtzv��mk�֘gP��E�	/�V��тJ2�䉉@?��1��|#VN��\b�k� <�(?��!�ډp�J&�m�sF�w8<��������MP�A��-��1H9#_OAsAʓz�n��l�a���K�/{��j���5�LM�F���=�Х4�X�1��N��r�k�=�u�iՒ�@E��M���ܺ���1��yķ�.�	)JFG�t~�z�~�R.�Uk�������Kz�g�����<fȵ_�g�m���}��ϫ��Z�8�z�j�l�>[�{�)��A�f�ž9%V� �h�1~����?0Τ����׶��~1N�>�Ͼ��4i�b�/ �B��%����ȡ)����W�/6U4�4-ׯx�y���@�_�ፘnG���+���g>������gZG�-��l�Lܯ�3%�B��6��p:��4�t�c�t}�1gL���3f�|��s�L���x?[<GQ<(1�d^4� ��m\���D"@ؘI�������W�w�j-�t�gK�Ga�R�1j�uh�������E�sG��Zo�ƌ�S~l�m��p��U!��������o�4���/�]����yh�W��ZDx1��}Z�F`ʓ���&pɒ�:�	!�$g��{�B��<���E?�3�����l�%Gۀs&ۑ�0y_`4/-i`������9¹���W����Ne��ݎ�NSID�����Y�d�����8�3�7�b��-�E��A��؎��O�;M�O	=�@���_�����l�ޑ��B`��w�`L�:.�Nꧨ�#9�E����J<ʕge ��/�����_��4�y���WN��I��5F��Uě׻�+,�O�-f�yV�=����*�G �SP��r�lϬQw�� �Oߒ6�4gz9�a�>����C�� ��KH�@�����Jc�k��ߪ� ��D����2��7W�H`1�q�S���R��-����`�'��M��[�F�z�����5]�᯻���w�����ެ<y�$�
fh�Nڋ�b���^���_�ͻ�u�#��T�N��j�;������ڦM^'AQ�
<e�FKS)���`j�Y[���=?��:E��;�w�,��QOu��GЇ=���8 c<����]��ł�6���yj�/�
�;�<~�x�H�&���"'�T�8��B�dxNi��ER�̋�U.b��t<�&<q�c�M	�PU(��h�3�=7)u��I�@���xF(��E�	�6�[]ƅ�L|7
'���;�`
�ek��	k?&������ޑe��ԭ&�'3��ep�_���\|�DOh�Y͖~2�:�9.�z���)�q��!��v�b���U߃a~O�?cz+l�ZP8Ώ~�~���W7����U~m���$�22�2�^�Ǡgc�\6SBY����B~�fH{b�K�AYS8�*��Rl5|��'��M���w@�WK̓T��@���	N��k��fRK���$���UT���q^�.2Tt�X���q�m�[l�?}�l��d<�s}� �4c(��@d�\�BͰ��O������n��L��D�e���#,��!��%	�T��N�yټ��E@�)1�G7��}?_�r9�3� ah���s�g�x�H�f�fϕ]dW�D�Zh��Q���ZX��*��RFQ����EHg`?3�d#�"`\�PH��I�yk+��[b�Eg�}}[f�;#������I�SD�=�j 3���+��_��&�����h�dcI�֞́q
X+�L���w�a��x�qt6�b�D<z�8� \�ΐ����%̩���Y�	ai>0��Y.���%�6�b4����E�\1$-�b��JaJ�Z�U��[Q��FU��{�3�6�SJ%I���́h4ν̅�S�4F��Y���ۍ��Zb�>�`K�c|�����*{�-���ǃ��ȶ��D�ه��Z���ԩ�$�M�c\���`�h+@�|d��&���������as�hV=3�����f�|!�<{7p*�-���ӓ�o&T���Өa��������(x�M2�~�֪_+(�^N ��[S���1 b�C#�l�/��������}����^B��Ns}nu�Bl���}���J� 	��:�!�U7=��2���y����*��y�t�!�|aa��P�u�@�F7��G[S�vp9BG;],�T��9�AW��%H na�����a��}��7T{��f�֫�����T�3��=��F�y:��JqZRl(A&�4�XQj�B ��B|�2´���
������wih4J�%d{�!*����r��"m�Y�q�]�Z�-T�؈���V  :T괩�Z�&�K�A������!�4k!\ ��BuR�$�w�ڎ���h�k��H���O�Sm�&��	��ɔg5m�1���F���\ᾅ��dJ��[@�,ާrA(��/+��S�~�!:z@c�@�	8�Mm����DOp�:;N&������F� Y�F��"jhaQ��%�yR0�zb��{8���!$/A�Z˜��\��\ێ�t�]�� =L�X�i����kY�I�
��Q"T �u{K�2����:���YS��]�<q��z��=j��EXt��en�?n_�B��yp=W��@pm��M������l��G6�q^W��W5coY�쬞���k��O�ŉ~jgN&T�����¦w���h���i(�����1`����mm��'�7�<��x�a�+bx�n��e�-�S�Q�X�j1���!B�b�E�nw�꬘'�@��(�fi9	ٷQJ?�}�j�����,��Ѿ0�L壩-�U�F����}�F4��m�������(���3f��1\����ȅ��͍���u5�x⼗fLe��jm�$xK��܏a`�92��A�qI����c�X�ڹ�AU�_鲆��b�d��q��Q��/�P3��T�ɪ�����v	��=���XЋ�
�OR3N�~���QuF�3�y�*qC&X�}���>_a�Y �0B��e��'0g�Η��y������TɸWȏӳ�a53�q<{'�9M�D!�nޟ4�G�f)�̣�w&�!���As� g5�.@�e"S������@rZ��*�/����	0B���K�"Ւ!�繽�ǯN�п��Nčdb�q����خA�(~ރ0�]������_�J��1���i�3y�F^�V
��Y�ˊ:.�?����:7��Hۼ��K�>�F�%��U��������k([�A�:N~Caö��?-��֏_�G5%�ζ6�2Ln��(��?���KS"�},�׉ʹ�s�����\�*i<��X�R��?��|�s8ە�o�;��O�3���K���sna�K5�P�Y]װ摠p��$�e�ђ	q�8ΨhW�H��yU��[�<�]5���cH�1�7��,fWG���O��a��E��`^�==&i��T.�˴����ritq����?F�.��1p���ƀ��jL�/c��w*~F�[�Ǵ9�6ޡ�P��o;MA)��D��xc��ԙ>u�Z�E���}�ir⼏�h}�x��A!/':ٙ�������Ek�l���DFc��P����S>���9�R$J�iV���S�-tx/���J��k�=��֥�������Y�kE�F�	�耫iv�Hd��PԂ�Ed*��f7��NS�z����,���CG�:�����ED�MUk�R�H�%�;�3�@�y �n�Y3*'�<{ۥڙ,�^&*��&�v񺅗዆�핹�񓂼M�2?��{�ߖyd�dǧ�����sԁzN�$4�uQ����p�}�E�准$�5�_G���X�U�'ݜb��s�)���i�8cX\���h��$�M�\-HOOu<R��g���4񳄷`+{Q6V~�b.�k
^���nFԊ��%��~��-߇a�v�4G�����5���MT~��Nh��j��G�<e�X�;���O➪����I�F3�Z� �MB�E��>�./�NH��MF�p�ƶw�����8q�����e:A������O����y���lsA�+�?T���ȸa"+��D��9���Z�>�;��.ή�=����AQޑ��OS�A������������I�d>8r9�P�hK��/a�
�&"#waf/�!�s4��|��������($Ë$�*�%{�<�j7�|��
街s�ש��~-:�����1ף-�i2٭F�N�<Ѻ%ʈY�v����ۜ�n�In}ԅ1Mv�ws]x�|O�*���X�	�Z��<ynQӠ?���"�V`S�c��"�����PE��r*93�`q=]ݨ��NK�̴����R9�si�y�7��Ć����c����{�,�ЗJ1����x?�诎�Z�j�{J�E�BREC�#�v�=����!�|y9�P]�~�׶�ɚNl6b�Θt����BPs�z��R0۞ |�@)xO�#�ؚl��cw*Rʟ�^�Ym
�u��}�$�V2���Fa��*�d�rvn"��w�&�ʃ-�i��9�o=qE(���~i0��H�0��[Y���T��c������
��O&bF���')5�_�����f��|�Z�N!�n�6b�ɏ����x�N_�gҖ)K���@yocT �&�tTw��}4����yȄO�y�a�f�y���Y�6��e.@_�X�bT����Ub���׾�O��j�w�A�<*$�!"���3S1��g� ]�r)�_��y{G��U�
�y�s�~!�w�զ���M�Pȶ�RI�k��5{�VM���8_�֎��:�Rn,ϗo���&�:���p�4��1���;5C��2�a���ȍ��}bsONQ�=�K�J#�cH	� ��k]9�����s�%��'��2,�s$�z�cR?Ǳ���H`Mԓ�{a�ILvOYܕ�I[�r{�Fy~���F��ot-��+��V��9ZYc�%���XPV�7۞�n*���А��.%�v8���t�s�9-�$���@����:�#��7�����nU�x(UZ؄�\��}@�y����o���Y&�|"�B���=�y8}=#4��\����f��9I+.	X�uT�LB��ê�:� �)\�̉{��љ�}�ߥnzh
DUގ�ggo��R���/!<�G\M���Y
���В���m�N���*S����f��Q�J���kт�nB!7.'�?���]�b�2T�o��K.��z����a�h�!��
L_⼅�I�׽Ik7�1$��O�IA�#6ݼ��U���A��=G1�哴_�ZD�%L|���}�>��;z�\����G���Z�R�2���zp]�PD=/���o��H<�>���5p۰����x��"f4�5^��G�*5�$w⥕�Rԧ�F��P����Oq݋�}��F<��W&����9�ٹN-L��c^�U=l��*��;��o�>����p2�p�k�V&�gG�;�4��;r;7��n�#X���}�ndJ�
��q�XV��W)�,#]�����0����X^���$i��m�����_S�/	n�ֳK������ގ�V�K!=I�PM�&qTF�ڨW�	�![�wX�Ȱ��ς�e�[q���Rq֦J��[�y\�Ҟ�	�)�xW१�	�4U'��*Du�����	�
�t�N����KC]M�ᷥܓ�
���1F���_�`ӡ8!�{&s�ט�է�d�L��������;� |1~���J���Df}�sq�����V���ߦ/����0I���s�Su��_%f�xN�F*�DG��: %�>����Q��k�	�<�߀H��+GW�>5iƒ_쳄Y>Eޛ⥃`@���@8�%��ﻄ�h��kgNJ�p�Ӎ�qT��3�d�~�։�ើ7�0����^qg�Y��o����q������$�ww�xi��Niѭ�5�N��
�y�h��D�
5�I,8��5rg�e�XWvo��3e�.g֑z=SXd��#̈́(k��P: Ǌ~6��j���������Ҵ��:�p�}c�����Ҝ�~�U�{����)����x���F}���P�&��3�����a�xeM���\c5Qm���9��W�^l�r�����a'� �|�+��"�4�/�q3C�&�q.ψ���.=��V�LhA�ܞ��S�:&�H��|h�W"J7�<Ú��mM-�<���n�oJ���N��[�u=q#����e")�kG[6J������,ߩ�������U����{>�8��0�i���h�+������?62>�����b�}�w�<= �ŵ%{o�7o��V��%r��t;�R�f�@r"�4�DG�
�+�2tDO	�S:;V��A:�c�����LI�P,�2Mz�������.�������z�ЩB��d<���mU$m��l��X�5� �=�2�$��6�P���Dzct����!�ͫ�O�3�If��\�d�z������T#_��+��v2�R/͇�슕8���:S���hf����"�B��6ٴ��Aي(R��d �P�`�;��)*8E�R1<D/dhy 3 �ï�6��bǽ�|j?`N�h
��O� �M�����s���tjs/�s��s�CO�5/��R�5v�96�D:Ϯ�bVY4D���U�E&G
�Ү�����T�%ˇ�lvW8Q�;A7��L�RIS��w�:@ 5^_�F�h�!��Nz@1)�U�a!�����򖚱�oVj1�-�O|	����q͍�D���8���!<����)YIjGӗ�Xj��%W[��U�=�.�����I��c�Y��[�E���W�w\�F�<HU�z48c��yD���h�Nѕ�����2�;��$�.�wU�� �V"��}�L���o_7E�(<����Ī�^�o@�p���@��m�z�G�P�Q�ŉk���l s�w�ۛtE�1p+�4�Y�����tJA���h��ie0�	�o7�R�����A��N.el������%��d-Z2:��y�&���(JL�m�Ѡơ���\h��J��=y�Ի�ک���؎�*(���|2��V�x��BT��pX�.vf����Y��-AU(�
�O_C*�0%<aj3%N'�(�)Z]�2�f3�[�x���ũЪ ���y����4&����������,Mɫ-O��#�/oyPm׎��ϮS��F�|ٻ҇0��ao�j��=������&d�<]�Eht���:�ɗТ%z]�c��G��$D��h�>V�
ծn�h�"����E���B�)6��t���ȭ7�2��?��
Y�;�z�c,��d�S
���g�X�}#��l���(����c'���YÒ�rӠ^�-|�`�PT��wF�����?~ ������_��`%)G�l�:�dCl[���#�1v�?��*�d�*��ܒ�D¤(��5�68<� �C�O�����"�'o:%��M(�Q�֐������f$����5L�٢��L� ��S1P]
���f�L�oVKw�\c��dF�vK���|��,Q���
���ǹ���j�C�r�_qz��(�5����CIc���%���B�,�|��\��,p�2s�ͫR9��P+��*�3�k�ꨄ���:�t0>�(^�Ŏ��0� �uq�����Y�v�(����F�T��Qݨq���g�/���qp������<����>���@�������ҹ�d�#�nT��� �6YV8Ԇw(�ջ��5�E<�k� ���&�F��NK7F-}��N�_X��o17�w���<5n �eS����Γ:;;�Oo.�3�����*�¨��%�AK��r����?����Q2珘��=�O<����w���Ć�@�o�+�D��d6~�Ҡ�b�.��6x��#׺;����|��hm��9bP&�����&� ��%/4��Z�&0>֠Yw����L�ozś®C&KR�G�%��z�r�5���ЬB�����r�"VN*���#��s1n���Z �s[:{�ki���(���ߪޱ�n��A>�&��+Џ��뗌�0�7�a�B�Êԍ*@��4�&�"T�`�d�K���N&� �yq���Y��)2�L'���#X_��K���*�f��U��76�֢<
O�bR�肩��89��u���Q[/��:Η��榨i��*D@%��� ��M}�ی`Y�y�-
���xY�Zy��UJ�=O7�fk�0:Y�\maS5��ʲK)��_�	�\�2H�;Ž�|;[��]�C/�l�U�o":w��=U�2���� �D�I ��]A���*R��;)燔gQtJ#�͌{ԡZ������Nj��"���:��na⃡hڒ�ԡ�����pt���u]	�z&����\1�]R������4�D4�A��
&m�|��b_HT.k���_�����puM�#^ypg��8�������)s1MG_�/?y**B_��e	��Kz��V�L���yG���ȥevzvkV���N�`���/e��'c��wyV�Q�ty1/����W!���M|���\~)���.��~�(a��������6^�/�f�Z��dd�F�ө�ԮE���[��$�R���P��k��b�^��.�g;��U�!{/oM�%m��[�ЭL.�����g�㠦D�VW����d�ےTv�&b]�X��������[��+d���im�k��< ���� ��|Y��8p
?Pţ{�Qv/ۤCΈ�쌬Zկ��"�݆�=�R��%`Ռ�+%{����n-����i��u����<�`~
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
���[p�Ky�-	J�@4o8���M��h�tDmA�c5�rC۠
� 4��/�rE�B�!t%s��E��@���[�?��M�x�*��y].�y���5���̝=3�18ǉ�7�Ȍ�א}f�$����ܗ��{(M%~��E0���0�j(z���~d�d�{c�ʉ��/��0�B��;��`u����KI?I ��p�Ԙ�p:�'�Oھ��Z���d����f�XZV�I���El!����pz��5�͟b�΢fe�	����9�/;��w��ET��#�Vt��}�u�SV.8k���sGR��T���֮.�����gF9$C��!K��v��C��o��G���ͮ`��J�����#��Hz���}���@`6�H|:�O����eSYV�f[d;�ab�e�"�Z���v~:��8 �x?e}$;�n��5������s�F;���R���^��#S+�csb�Vi�8�+�V=
�p/!/�bA���@!�+g�<���R޸%����<�K�[TxcUD&�o �o���#誦�b�8��i=���4� [��&�V@��k�aÃ�~�Nɜ�^�N��\��O��a8��6��7&�����˸%����堎��� ^���H��&�WY�B��?SP��+��ӁYzꤠ��r�_�ǣD��$�W#̍��H"�����\;�<g�~�s���v�w����\-�I�ǽ�|��w�[��@uѸ�-�ɉ_B��^�"?~�`�ڹ�H9���*~��!r'���ܕS��7������wW��8�s���J�@)f}�Y"b\T�`GB$[�L���J}g�������������V(�0��G�fm��s��f ȲLc���Ӻm��]Oy�{eݯ�/V������8�m"�b���Os�G�縳�P��W�kQo�R#[�ʫ�P�|�)�t�7�p���ݺY����ȡ+��3����s��ɖ'\��	%A0"��ס0��nХ)q���{,e�U ��;��i�=�fp�g&�?qC̬����)���v,�3���b���(�Z���o�J�W�\� )��1q��ʅ��߆D��r��wSM�4�v}��b�M��o��a�%�Lbh��d�%X������B���Ja'ݮ�: ��6ɚ��Y�n��FWS����U݈�D����с�aL��3q�S��u7�ec^��u0=���J-�e���ŏ��0�4�ݥ�K�z�$o���e�_u��u���.��o���h�C�W����R�2�U[������h����j����k�F'��]�r8á)k�19z�sɬ�ٝ����}�?��(��{��!K�8����OI�Em��75��$�����
Xr�HQ{�L9�AFW���dۆ&�a���qA��p�}$vu��Okg�y���.,���w�8�z��%oLɤ��x�2���u�oUe�(R�줼�	J�w4%�Zf=v�������{�޹S������̖V��t�5�����̭�;��InL��\T�}�Z *��;g[��x7�MM�o���a�5��ܶ�}l#��'3��&G�� $��f�x�q����[�ۡ� F2��B�N�߯d8��@�|=]ni�:9j;7]��v��L�u�:�w���Q*��xt�᤟��c_E�+Ӝ�#�f��}ޞⳚ�p��c	���~b 8�%N�M�?M����6}���XЋ��!�|MTh�&�M^abu/Q���~��(@��'�]��ж�_;B�I�"y�z�GI���������_�|鸯���̖��}S��=^���|�����8�Qj���[s�t-'L��S�+�_KQPlakue�En2tx�Pw劖[�H�7(?N�'�׆L�f�b�O������=Q9_��`����-n���~Q��&�_�,�z�O	��k������h+_�Bj_Jﱴ�o�������\i�}��j���8�΄~L���5�{�5k��r"��$��l�i2WL���a^��d-]�1�r��7+��R�\[q_��}6���gv2+L��Q�-~�v�g�֬�_���ȕ'��<O�y��@}kX��U��{ڢ�9�N���Lr�
eNNp�r��g����g�ū�{ɇ�3L�&D8�R�|M���Ri�/��-b�jU�.���ɏ)�̧��P�`�}ͷ>�|�Sue屏�&x[1�h�����e]����nR�Ռ���}z�@wbd����z��\��uuB9�C�j�w3Cw�_Y����HC�= �Ry�kۓ�4~z��_a�T�o��lQ>m���B�цV�S8�{�7�v�<O%+�D{$z*A��&9��u�WJ���Dd�<����	�F��O�׵OC��h#���ƅ�A1֍��w��P7���A�xkM0����}}:+e����cm8�\�>eq�\2S6���M~�i�S9�4�)��P,̜�ش�Uq����ցf$/�<����#��I��c�q_d|u���=t~�Z�n��p�k�ۢ���$��;��a�Z㙎v`�F�V΢Y��d8����%ǉ�'���v߭��e<�ldYh���F����7��ϊ�*g�H@V8�3]/�n4�������
?̟Cz�"����R?.U�����@��ܚ����	�X>WA�:��W<�}���p=9Z�69N�V�tq�����~*�0�Z�����T�[(t��F#.�ߒH]{(.��T�S�ۃ �4^ ��دK �u ��mb�0�3��Y��C�`u�����]�]��|���FN��\_��(R�+��`�w���	l&�N�	�!!�1>>�2(���^x����A��6-�m��X�K`XױAE*X��*ԥ��ye�B6�)΄�9�`I��^����1�H�?Z�+��q�+��*��nH��R��͋���0�#V͋w�V�_��h�w�Q]Am.Q�4Zd�#���Tꃐ��7N��.���WC$݉|$�q���I��~��RX����뀱�^Cd����v2-X�c����\�QH�14����M{%�Z1�}�y1G���Og��}�K�S�ޫ�q����}��.Y�s��,QQ��qb�$_+x���
��/�T�:���l/�-j`�u��ڵq��k^��
���BN�]g-IU�i��ʿ���=�[��*&t��Dt�QV�'���.�ʭ��a�vo��-��얢!RF���H�9�F�ʅ	�ؕ��T�);A5�r�����7%�~L�4���?_x&O�(�,9z�ŬLr@��P�0=��r����尸g���y#�x����UONK6�=DӮ
z4��*F�ж���m���ɂ\|ph�{�e�2�OfT\q%�3Ժ]�E��B�������2:P0ȭ�(�T����;	�	�ƑB덪$*�#�!�8"�k��A ^G=k�r�������m���@xsf�+>���p�+ם0����%&�a��+��D�&� �?Z
��qEƞK#�Y�3�����m�\]})�%��BT�D��"���8���1����E��2���CYD\�F4���'1n�����c,=��4�rTT�-�{�!	�"c�����)Uy`������}��Zv]�@x�������ᕾRsH!���'e-K��F�[��/�N� }E:9�(&Pd8��_������� ��$��F�Vk�tw\��������/$�3��|Y�/����K�')�G�"��ִ�>�K����g�h�S�Pa��<�Ϣ�."�#p�l({�� �2���ꢖ�.ү#�(S��+��S� � m����O0����2�q�t�X�!�xJ�"����)�&M�+;�2!��(���_�7�J�߳� g6�����<+1y.v0��yy-c�<��U�W�8�ax�a��?�2G횠���X�?����ي?��n����R�����h-�g�D�-��9/�F��,�`N���il{d�g�#��ޒ�Ed@}rk�; �+�[����):/a4N�ږ~�e���!%�9Źj�K>Dm�e�ѻ`�Id�� �]�H�R�����I)�"��o�$(���g2�m�@; ǎĻ�:|�.wjWSNj9��"P�ۛ���������t�Ӕ F�>I*�p���	lQ;�H,�uu�B/��*x=EM���B�n���Ⓑ����m�&��-"A0ZV��!Υ��d�|r�?}�!Q�%�vV[�����(�K2��q�<�^���t�k�����a/��d!u��;G}�4�g	�x����x6w�F�vrJc|^r�E�|
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�
#�i�MS��Q�
<B
�t?{�^�z����$�����Yp�Z	��O@�/iO۸�3�����p�`��#���+�B�&��Tf�O�}�li��x������2��c$����<Ԡ'��Hb&�[�q8غAC
f������8��]vʝu����@���-@�0{o>����;��9���1!(�g���?�
C9
e�Y�[� y���Ts���b��Qu
�;τMk9'i�=���h���\='��c��+����墍�n:<��UN0��k��<j�[�ȋ#+a�ݨ���Y�z�cc�PK�22L��e���%��&#�.�Vd�Խ64ʥ���w��aL3�Q6�t�*~v��P"SuW�}0~3���7��0&�r!��\Aul|���b�Y��th����|j����i�i�2L�i�p'�����K)��y1��Y��u�ȭF��&�-�:;6A&���7����nNBj�Ho���H���?r�������݃�&˾�\��2���X�w�B�25�n�<�����Pc��n��u�M��xCOK=�+��Y7N��N��d���]���Ȕ΁��h|Ĭs���1�7�z�N�ٙL��QA;��A�1	2X!�������n���Ċ[��TS��e#���G���[�13Y��c�Z��Y�TNQ-�����I�{B�o���Q/�kdW��ϯ��k�\�N��n��as㲰�J�*�I�`��vk��9*��׭�a������΀d)�_�~���W�C8���t�-���o�J� �煾�xbߎ�/�&�-8X�����,RW ����b]�--c�1�4t���7Ќ�4ׄ*���.a7͖�HA�4H��o����~��*uX/kp����!��O�,{9�Մ"Y��F'l	6��;@�WzB���{p�8�jl�8%P}��8
^�	�cR�7��BC5�0��o3�!��b��͵��4"�\[Z�|y!��� �:��}�¾�`7��^[o �3�Ss�(�� �R��V����q�C�6σP�z�r{�U��퓒ᔴR�-�v��Naf�u[m	��´ŧRέ�:2�#�N�
j�0�Z��g�������lv���uݝ������KΙ?JQyUvc��5i�)a�����S���HYML*5_#��Eo���GXgC�I�*[45���j��n>wxA��fNZ��ys�7M�;AqC�����"%�5)�8Ǜ���o���u��h�8A���9���m��Li[�U�u�lߍ�;+�#�!K�[�h���'<��N�<_���ΘB|��}h�jT$���	���R%�Zg�U.�lJ�9�k���_ç#�Z���{���:�B���t8xoY7���2W�"6��c���P�)m�]�_y�#9V�oA�{7 ���K�םT�d.� 7�y#j.X�%���$-�{��Q:ߓJJ͵�����Ȗ��/�p��S���}k�:��Y��[٣�9���<s�*���K^�0n����^f%���A��D�ݲ���yǢ�>�:�lu����� W�j!e�!�`g����B��q�E���Z�J�ެ4 �h&&���4�/q6����X�t��fOQ��c�4�ΐ��1��(�a3�ni��(��h�O�򜫓K ����Y��e3O�کg7�J�9u(o�MV�j��5���p^��-
��3��N��PIծ���.��<�@���{?�mlJ���K����R�K=컲�#��꟢+?c�y�����C@�+M�s8��^�}��C�������VV(��؀]@>�'p��(փ!�mh�#��ALFy��ؕ���*�B�.�D���cr0��"�𛋥|u�=�>��(E��ޱh���!6���=[��a�T���
DT�j�q��ݛc����I��3F�׏@D�ߟ�}��1_ǥ�̝�/l��'Hb�8E����1.,䣐J�bc%�	�)��k�
h<�>jn��%�-��E\o+�&���O����9�~ʍI~u:��=���\�;T�>��"������)5����s�ζ��2�����ʈ<�V���6�$e�U�튖�#p��-�c��$��Q��y���4,b�Z�\�\Q��]O~�N%O�;��s�[s�$���D�I)M���#��g����~�������S_71a�����Bŭ����ɭ�v n�������������Q�}�)�o}�_��bh;Ӱվ$�V��G�0T:sS>6���ϫ��𞱙bSq�t^a=?������5�:7|V���m��R��=�K�<6�����90�q?��6/�<�lKU2���'�H.�D0z�t#�R+K)�.����]�>qn�3�v�"icqFj�%-u�!炦}��4x���[,1��y|��0��K��;sőu��D��*4��3�@���m�hKG�����tH~�8e��A/^�p��l�^C(�M�̋gF�o��S�a��D�/�ǌ�f�3�'@#��$�@��\�?�CR�x�1�FYĂPb������ �/bܓ�X��u�{8�t��r��;�f�JX�!��Bߐj�m3Y!���(�!�*�� � �Y�ο�ȝ��@ݲ:� 1�D����g�$��%�I��J'�s��;$��w��"#��!-J(2,4�q�Ԙ#�6��K�b~/f�xj�X�d�l꣮/ox� �����m�w�T����e䛸JhA,�c���L�(B�Gɖ�!	��}��OA^�qH��@�ɺƶ��e��3^�+l�=�'��wU���a��6��m���XZF�Vˏ�D�������HK�� �^�ג`��� �H����������O�" U�G)�f���c z�l���޳��o5!m3�<
��L�3=x�7T�򻶦��W���:�)br.l����=>
?�_`��зֵ�¼��!���_�ш/#��o��Ϻ�h�~$���B:������A*���bq��u�K�L@��(�@u;�	�n���;X�HKGG>3���%ݫ�?��R\ >;�V�ɩ�����%��e�Gѿ�׌� ��je��%��2�x�w�ݘ��.��xӊG��4�s#�Ֆ�i �
��qH���ɏF�7�z���Q���$ O��9"5�U����R��62��f�ٍ��������X,�'Z]�n4���
g2�c	�~�)ü��Ha�G���|Tj��K���A���!~/	�nP����o#�0"qĨ3�%�p?;���q�����̹ߓ��At3/X�Api8���Y����E�@s��;'�s |�@ m���(v����tt�����|��w�9�mUg1���	U4cl��`P�¯����Q���KE�Oj��v�������J��v8ohtA;H�]�����k#��7#{9�a}�$�����i7��!�հo湳��}��2w�߇��}�X{�nm�̝�W�C���������]]�^c� �/v��=X}�i�[U��<���`�2D��1GTj7¶QR$���*Gh�DXZB���U��i�5�B��`�P�8�j�nv,ƴ��R�	0�Ou)�4MV���Y,2����֝�E�a����X�jr,h�qŔAc�@�9��gV+�ʧ�,�82E;� ��2�;�bU��U�����+4��-��������2���Ӳ��g�(�e�j*7I��	����I�g���^��*׼�7o��&�\^#1�oI� J�+Nq�R��e��!#@��+ݮ=�X���s��"Q�����K�r.�+<��c���
��!����"���6�a�=-�?+��Oz {�&cU��`d�ź��F�6y�^����h��6��ot�f9H��'�������)��=��_�4��f.+^m�\����}+��Mnw-vI��%@��];�� !���L�s"ޘ��;K�6�^KPjι������SD�6��@ߝ%d6�}��>Y��v����r{��i�&Ǧ4n\�!Q���49�\���(�ŕ�4iC���	�I�@A����t�L�0�QG�#����@���r���z�nQ����j�/VH�D�[ ��8pgEA�T���f�"$!��AO�vY_Q�x5���7[0�zT�'�p��#�f��ia��а6������:�y!)�<�WdS��u����`�ꄌ���t��nO=��O��L��+A.����E���e�)&��YT͆N��Ù���d�/�G�P��X,�0�ж,7�#*u����Y�a��h�C�%���5$�ML��qFBv�ŝn��<��]��k�yl�Ȉ�.X���X��JV��%�l��Ù�9��$<�i(7��Ta__]p½.k�(Zn��3�+U. �n�Z�nkV0y��˦��!W��I��TD�6���>�D�> z�9���Ą�w�u�.����Q�c�ܷ���l@�W�7����(�!�3yR��M�0�b��W�ܕq@4�G��g��g ֫��;��w��L�����%v��qmF����Ea!����.�Ώ��{��ϳ�����D �#\���t"��i���0}��Nqr�IȾY�#�#��`����4����?0�����c�e�Y#&��+�����`��Ͽ]v�	�)��O~Q�����y͟t�]Ɖ���q�:��N!�Y�2D|N����G7O:��3:��e�0�}�S�_5y��џ��ul���Fė� a����]LM��bO������;�R�$�z1�7�\U��B��Б���p�3SK��+���}@�5)���� 3���`t�cLo@�9�#h�kz��^��7�ů�9�/�O����yǍ�>p�����AP}z&�A ��ѥ8�	�C����|����b�,���yD�3��fn�U]Xuˍ$A[�:�}t���y�����U�=��CA�o����
��p<�}Lkv:���{�w���|���Y�����S���Dxp�2Gf�:]��K hO]�)�MhL/���[�h����K4�eg��N�(��{)� �O�9j��� �~ƪ~gh��W�7Ok׿�<XP.��ȴ��Mm��)�/�.�����c��!�W+MZ�4q�ɵnch��,��ZJ� �SHE�r+����n���`	ҿ�k#8cv߀��n�� ���c� ������[�6M
L��uVy֫mŮ��'�A<���D���e�E���"�Ч����2 �/Wf�fLΰ�N\4Q.��?���9_-�/�
oLka����)�f�H�O �.��X�p�#'����Ӥ����)#1�;�}����8�Ԝ��A�6OV�MD���L{��ϋ�As-9�	��<яdF��
�o��9����LJ��aZ�O8Ǵ��7Y�����a��k1I
��b�7�%�h|���Q0CS�K�;�K���qFKՌ������)̕B��jA��(��@h^�{��G;V�X�xϵ2��5�������y�R	#D�#Db�r��E.B
4i�^��4����A��$�����WP ����˥*d��uJ��8ړ��(T"z.��:CD0�V��9����+΁���)���#w8��x���#�T�V:�����
��|��b����{��E�:�B-V�vVui�����Q�.����S�
�	y���?&:rȗ���&t��f�'����l�aR��%���ڒ�u,�Ѩ���1h���@�21����]��B�����7�F������~�.�tydCG�9zG���'�1�����*ɺw;r�e&�������B��M�����]��_���*�M8��ߝ��9/'mB�M�$��)��XK��L�0
�F���3��֌������]B�}�I.^�Sbڳ�]
�)Oxp�P[=;�I��`��������1H6o�d�Wb�㌲�ňְ�)!̦�w_<��p>s�z�p�1
��ٯR�?�F���Ҳ�:6ޜ�RIV,�������U��nN*��$K�F����ϋ��I�;�%�w+^[����Y�{P�>c	�Lz�����P!+v����m�8n��;b�v7p���|��u�_��A_�N�9�&��b�<�E��Hr��ǈK(C8����0�#G�tiEH�� �H�9Xc��Ni�=b&��3�^"�w�xӸ;�ۢ�5���u���<�mA�m�%3p�1�� �[5�n�r��g-�u���8�)z�N~h��u�IM_�7���5���$Vb�9g�/�&qai��R����IB�a�t������Z^�������aq��u�=��yA��s��ty��a)����;�I���L7aw妒?��e�K�]��:F����ߍ_þS/�,C�$�̦��qJ��VH�Ԅ��M(�ؾ��s��r�ѩ�O��aF�5fQ|βd`r�e6��pD���L�������e}�ŗ�C`��z������=�Sl�M��T^�����IjxV2��ד���^d�`!]�Ć�Pu�*8����{j05c���g_qd*}v�y�$�������ۈ���l�rq�|��j4�OUD
Z�H�Q-�ّ�H�!�y?�v/)������2$-~��!D%��1;q�ղ��!=腵!)���7vWz�ĪM"���Ԋ�mq�(����X�!9,.�nN�N�:����-��P3�y���f"mt��
|�x� kD� /��(�_��z�������N�,''1��H�_W�\�OY{�{L:\�6SmYЍ>�!���r����X�2�|�P�pX�JnC\�XRxuc�/Y.�δ�P�~��� �>o�U��&}��VI,��eXM��$p�;LQI^ɸ�8Io�i�'�?�[���Ֆ}��M-M[g���8@" ��	>����ϴI<�����k�Qu�M����犕C�=�{�P���ӽy$hb�ŝ�Ȝ>x`�7���8]q\�)I�W3FX�!�	X�����x�S���c)�d��A�f��$\���4b/@��V	�k�/�~��ʪѱ��٥��K���cȌ!@U���y�į�C@Ab���S��k�<���˵���V!˫�([1�a�>䪍���y$	�oq� ���*�Yl�L��Bo�,���
��6w��N7Mq�&����a~7�R,�u�F2��4������[���lE��4d�ui"�=��{�	5nIwL&c&��YS�A'0r���P/�?����RQiJK��.����1��X�.)ER�x�oҝ��0{,㻚U��"����>���{a�I����
J��L��'�ְЦ� �&����eM��T���:	��C�I�N�pMU��99�r��`��ͨ�YV߿�h���#d��~��٘6�/rژ�|�, yqHWO����Y�W:�9,�R̀}��T����*�{��7%���刭4 �GZb��\a�3 0]���6��<�ڭ/v��_���ڞF�Ln��f`�!y���v�d�Kˤ���:�I��2�g(|�P7��{>\%*V*ΐ����{�:8K���$m�q��� �`k�I��kW9O�c�@�Q������dĊ�{�V�.��&
��EnűBy�L��V�P��B��7�`7���+ c9������y��]A�Ƙ�B�Ҝ/��"�DFM �e�ٔJo��L1�hZF`�jiHo2���^������"nT�J`��)�I�T?�[=�o�gHD`�E]ih�|X͝Pƅ�p�Y�rF����y\
rɗOs,��%�̀���|�C!��ߡ���]��h�ΖAkBO�����Y��j�mC�N�z���1c	��*�ǔ�v+�w���/e_���������gbB�Sɍ�lM���Y}:�8D�1GH���fו���º�P+z���|��;��hef�}���(����Di"#ƥܘ2���`��A�,����2'�ArH�hd**)��+��j�,F�l�{淓'?��.Ί���&�Osrfx05�H,M˗s�6������z�������J�.���"?D���\IտBA��>�����F�.-YMZr�O<��X�G-@N|��� ���B>2� ���b�?B�	����e]�c	?�4ñ�KB"G�1���9� j��p�����U���J�BB^5�?�nD;�RVG!Xw��+ik5].����AD��/e�Jvg��$�}��4)��	��E����T���Z��FMOH�z�-��~|)-A�.,`K�N/f؍�@#�@Q�]w�(�1̫=	������QXTW"�=����*���ܱ�������'���iBao�.�<wc@�Y�"�:V���vǃ��1ҙ2�׬�����[�`�>:��~�V�m,a��P�0����I���s����g�k��oI`=n�M��4�9(d�Z�ײ�[mt/ޟ�p�ҧ��Ox�pb&��T��8��ɰ��*�[�ڷ�݋=�D�+ꢍR��h�g�n��ޱEKWP{��%����q�`�#0j4�'ڈIx��?��*֝�0��ugt�n֍H�t�
������"�?Y<I�qU����ˈ�q�����q��|(~9�I�z�[��\���{��-j�R�=}�jkظz�g�l?���U%G��u���9�8�r֛L,�����̇�@����ч��)�R��2u%��ˤ���?�%��Ò*S���*��jq��nӷ��S�{��K��Ғ��C;
Mc8�	�9�6����'G��;����(ڝ�BX�7*�~�Vd�h������.�qD7�Ƽ�i�h�γ���ֿH��ä������Ƭ����e8G�N��KȯQ�D���>�[ic���xN"d--���X��JX�Aߥ8�ڭ�.޳�*�-�z�dZ�u����F{M�֮W=�����K�Ԃx�˖���x�A�<+�0��Phf�*]{���)�@��2C�җ�BӜw�ٲ뤧[Tu,�(�U��C����hʋ�'/��Ps��=�JJ��8-.IX��L�[�S��F�� �]P��P�YȾ����`{��^ҽ��y՟9H�FS�z7eD�[)���i�)����$l������S�-��(T1>+</����ip��Tի��8�ߡְH�-��`�bm'8چ��F^[�v|��sZ�����6��𿟃��#Y�B�7ٸE�M�u�Z��/��xJ��O/���*.�k�<�g-����迻Zߝ:R'sNQ[]��+q4�»�7�92���w��Ѭ�;z�������'�nʏ�u�������ə��b���W��cܸ�!_��+��&? sM+H	���?I��q�!�L��_����N�`�
m�n
W���Om3^��>��S�����G���� �m���~0�d��FT�� ��Fb4�U��;��%�c	O�������0�bΣץ[�է$�dgv�b-Z^���5�ABSMTn���Qܥp�>�T Ӷf7�ڞz�^����a���R3	��@�Q�$�B,j�H:��ا1ȝM~�υ�JNe�o���U/�VHs�T���Fj��XeW�;�j��=e,}�b<3�J%��	�Y���q�-��w��!��m>%�,'���&�[ܑ��ħ|�2x�/ܹ5�ƀt��<��Ck#����cP�,��HCX8E5��a�[�5�BⶢK��Y<	�9���{�B؄I�	'uL�umlFDv���f��{�
 	1e���.߽����ڹ藀'ܸ��P�O�<�|������!�2F�/RE=cEm�-������:��/�ݾJ�r��J��D(�(Qͽ"K�b"Xb,`w)����*ή��-�ۡG�[>�B���
D��Gy� ��D�XD4.��U�ah�K3aϚ��v bz^�p�Q""bG%�n�{h�+7߶����n��-�g�2_;ۇ�e�+HR����Q��^6�Ѳb�M�ee�r�P����P>	ua�m��=|���1�h�H} �>X%�C_G��R��;�5���������ݻ�\�z���ۿ,���M�sz"$�¦d�kQ��虚�B7>	}�P#:�0����G�u�7�Sa��'���9|{	�Y�����C�f��;�[�k>{�)5�5W�ك�VC"�ݔLO�@p(����9���R�+�j���%J>�⒃g	�_�C�1����s2���l�6���^W�մ���2a�֟wW�D�4������}%�:�$`�9�d���n�{�ĝ��z�no �_���w]U��y��q��%���rF���T%�����O��\�%��u�R�E�5}>�w�?�� �Ȩ]�(�I��ۊ ��u�i���w�=��į.���<���ٓ��:t�x��怿�'6!79�E}|ʀ�^Ƙ�,O��~���h��]e�`N���
X��+3*�޼��2a5��s0{TG-7Ƭ�D.�'�ę_
@��м=��=�����ee���z##&þ�ıGr:T#�$Ɩ`=��������;�ifV+�D�ӤgJ��:x���l��"��(\�������"�K�0Ύ���&���,�c��Mo�H6ԗ���H����Zl������0]��=GXG,�W���b�/��ճ#tlJ4s��>�o`�tF�Tj������	۫���-�U��a��3�wIA�&g��uC%��{W�V�wv�Μ��ƿ��OO�z��۟f��}�Ԩ������~P(ZM%N��� �Rv�8j�fa#�7t�H�&7yrz��Y*�4�2i����B�.�����1���O@�	%9F�$�l�����j�D�o}�5�{ljJ�=���_:u�\���s��_�b����/,u-_@��A���X#�y��X��)I�d���m��i*&18_�T$z��ь%���<M����㪠��@��;�s�����0��3�q2�#�2�dw��F�G��}�	�����^��v+�%<]�)�^}.�+R����Ch:�^��bngr��욢��}�2"[z�ђ���h�N�����~�튜Sw��dn�����
�9��-CK`,�X�	��1,]��y�����.�n���>&w4�c?0��1_�pA�W��hS�����ǖB2����}nj{"
]���-AoEj׀ ߵv"r��H�(�>;���vnk���K�n�-s��t�a��oЄ)�%�S:��5l�w<��V�s�j%�U��K�z�R[�Ä��%c��d�M�������Ƴ4�r*�iԚ��o4��a6L�L�ʂ_��u�PRI�	���Ɖ����\&>(�P��>V/���GL͍���P��7j[���A}	��v%�x��#����j.j���rObHYd�o�-m+J���,�)}#2��#dZ��T$�t�;�F��؅v�O��?��ԴW����x�T����d����_6�eW��FM�-s�[5�eI4�Y�������������h����Bmŀ�hN�nǦtĹQ��.�˱�H��@:(�u��	h�@Dk�s�
�m�e�Z���q��A����5l��w�����M*@{ԧ���.w���"��tF�v�����hA�տB	k�jf�(�PN�sr��6���lf:���Z��$U0
��9C/��=F��F�����Zu:���wV��{ZYv�>��9Za995��_�P?e}Ȅ҉Z��JApn8O\82�3��
Z����@�D�2j�1�(�����Ib�%�#U��#Tk��k�9Wh����Y�33*���}��ܝ�coc<���_�I��F�A�x�D8�(5��'A1��F�
�_rΊs��ɂcp�՛8*v��7���?]ټ�kY�cSex���z�{:��a�A�jM|��#�y�B<b*������Cߩ	�oazÜ���� k�w��y@ldm�W�I1A���4_���2djb��, cӖ�����=�;����Q��kl�τ4�u�Uu	�0N�P�~�1FT����9����K�dC���룰�ҶKӑ7�?w�8�����$6p�]��l�EP�Ea���Ԩ&�� �f�w2��g	�Eg#%<e�MʚOx�H&�{��OI�|.�`-��Q�%~��Q�TV�m!M(�r��p����+5/W�n=&��z�Ay����*a�i��]�9n��>���1�~IyB�t�����RX��z��I��	��d"�=�+�z;��e��h*���c�;���vPgVbz��YI��]�r}U�s�I���?�y|/��ܬ�{��J��":�|��
���O ^ѩUT>2?�eG���A�����әLP���6泠�0?:Us�>�
罠��d��Ed�����b�W�^\կo�!� 9r2�p������b�H,c�Lt�=��k5��-��NR~DA6j����k�)JƯ�J�θ��>��eU��Y��0o&Q[V8����.��������F�Q2Zl0믱��mH�PrI]�D��T�G��!YD��s���jD��A�c�\?��"@��)�o���
�]�5��W�(U{r`o�ĥ��YG��:����lz��Y����"�7�A<��/K�Ñ*p�!���Hf k� �x#065���0�Ȼ�R>�d���z^ ���́���q�^՛��~�	k���F�uyK�=s���_2ƼgVb	�LJ��h�s��ȁ@q�@�/�4�_���^wڒ��`�������߾2o�	���#�H�E���s&Ϙ5R �{��P���<��,�
-/_�r��8l�̓���d��	�݇�k3"V�˖���`4����7dn`c��� �A��(�Ǜ���}�G�4蕧����@k��VTW��� ����?7fh�/�K�ź�٤��}E���Ԑ\~�;v��XE8LLB����䵞~P��zC�
�^5��Ɯh�ORD��O߱��J�E��B0��u��G��d�ے0�~���$xn[q���`z�O��\�[R8Jo��J^�T%(b]b5��(�%<U����k9�s�ޤ-�'����F�]��cUl�JV�������px߰x�[��ؤa5��ަ�5d��Tx,ua�v5$���[���v����ߞ��p�$���#�����v��\S	�'GY�Vi�/�}�N�	��)���|�p�R���� �6�?���cK(�L���<����YL��;�� �1�cT�ݬ����Q@��#ؘ$=��߯��)�-À_��'[���3p[��j��Uɔ�b�g�����-;cȕ=��*��iŜ�������D|3�^e54�K{l0ɠ˫�`M��(���A��kbY�'D��oק�hiA�eS�`n����>�p�X�ᵈ�cI]�r����w.`r�݆�E�1��xd���[ܪ@�KҰE1����UX��e��3�����*�#���7N����!]r��
��T��[Lǰ�C�Ŀ�ڛZ��&C�LM?���{�Q��΃_ O���-2�٬>��|PlU0���+k���@a����MKN�tC��Я��hbqI�<�1O��?�]��j(�Y��L�E�O�ܼKG�XI�o�G���}���c"�{�!����_��[���`=�n���'�;=�D���u �qS��lk�6�O� G�ۃ�@��%b�T�ҷ��?��]�k�R��/���I��L�G19�t5X2���%���N��l�:1埠�n�Ͷt��χ֨�y_z3Ǘ p��R�R�V%7H�Z��rެj`=��"`��沸U������k�:|\<�^8#�rU��k�JB��:�����痢x�@���"s�"W/�X/Uo�!�~>�@��y��k�;�Mڑ���MV�1L�m�{C/��RЛ�g^���f��ji��Պ�K��qg���7�%��Y���6@�F @�����]�a�B�J����s�ִ�"&Ӎi�x/�f��e��k�7p,��%�2��u�Ֆ��̾ׄ�E�k�QI���f�χ���O��B�i�p{�W��s��`��h��M�<Б-�^�"�yT絇T=�Xw�k��nN����2�]w)	̪�~�x~�qnR��b�=�B�<��I��F���`���c")JF˺ӱ���I}�{�a19*{9_��/����dG�O;;�f�g�x��G�D�Ѩ�f��l���������hU�<xVzp=~��ޗ��e�����'2)/��5Iwqy�X�0˅���d�.Zn	���ja�auA�JL�:׫A��?r�@���:��=�毷)6D�йv��C��SԈ� ^�h��a�5�����
IoT� ��]M��z�	�>,E��6gc�<G"�>П���U��^I��\�ػ����v�0�Y�QH�I�����B��G����%���{%Vfcm⹔4��5��E���2B�z0ͅ3��U�DcZ��_p Wa%4#kV��m��?��������u5T�L�T�l�ծXN��W���6�J���.W�<���-��Î�M�)�UV���隐��<0�kU��6l���֘G�Ӧn/���h�m̐XV�`�/�(�V_�ۘZ����fo|��w������:����9����#!��K�=��q
o�o�YᾊX��yg6ܨ�ƀ�#CD���LΘ��ó���)gB.��m<'�3V�PA��<�`8[n��-@_�a�+PWp9d�%�[�~���҃8Ue���]�1"*6#.���C�s�A�D_�sl��J�C���$c
B����[�_ʐ�b��D�\/D.�a��k[�Qw�SZW���ea���/�b�ZG�6-�%\/��
�/����.��_��K���2�R��?O׾tP�'���(Fc���ϕ�7m�+~�(�����=����Uf��۬ &��Bk/o3��Cܥ����|ױ��4p%�/k��I��Uؗ�dl����Y�P��1d:#�Fz�1H��q��k[]V��V���.�����X��|QL��.�o�,�v��
�����Pu�貿[��D�f�&PU9"S�v̨R2��	�	�E�8����>h��v��"��uv�Sb�"5V�ק�j|��纼6�oP��g6����x��ڷ���	"e���Z�̰���@�DC�@��4���X�>��U?���ۜ4���ow.Xdʸ�e��noKD<�Z�L�l�$f�kn��4m��+a���Y拂*�\p��8�I�܏6U� j�gדaP���2Q��]����B"��0��_�����s�r�U����P/n�]x-����������0��b��k4���6o�p�a��1�HW���x ���8YŴ�rqd
�hyȀ�urMowKS�m�k!�ݱίK��s�N���JB�=�����'�<������I���s4����T�·t�)�Q̚0�r%'/�?��u�߿b�z�  *[&����7���5?@���k��J)h�1�2��\��-��_�ަ[���ϊKA�pny,'�&Cm�Y�qD$��c�+���ȑ�r*�78��Q�����M6=��
`�tl�I.��qO��mI�<� @�(}�7}�٘�,b�7<���W�@*^�Ѹp�_�r2�[���]��LvL_m���S�����1��;7�:-��U��P�	4^�v��^T���dn|Gw�&8T��F���u`~�r"���E��\����!�Ӧ�y��p~�����=yY+�����E�o��1��Ό���bi�sSz�a�o߶m�x<�)C��2��Z����B��c��5��%¯��1T6[�Ao_�<��}Ͱ)	�z�N��V��b���lDjyX3�4*�t�L�ү}Qw�}����k9�&�$�N�џ��CNVl�ui��ԟ�������M�̯��>�:::���pN������� e�6��yM��xR��"G�}��	��D��1O�w�3��Qـ�]aꊔ���@�~���pؿ�ls�H���)0�mq,(>����{G
&<c�q�z�T!_�̓=�e��a�{�ະ���m
����960I���"-��\�"��G9�E~u��U�	�H���-�l�I�z3�m�XP�D���6�9�%>�W�O��1� �[�8�K�C'��t��P�n�����4����,a�ɷ����=b����ע��xz��v
�)�i��u���V�c��W>�b7~+��o�K�ڥ��ӕ.���p�9���v�$��]��yq��t��G������v��l�����W�=2#|(-$�_=VN�����}���c2j�N;��O���S��(Eۋ�6���d*bB�_ɱeڲ^�΁�d*Mc����v�@ ��Bܾw*�GTS���8���RM��n���ί�+�Q��}��0�S q����ޮ���p��a��Gy�!�]ښ.��P����E�����֗�]�O��w�?�����(,;܀�]��T���~ɣA�T �Lo�|yhMz���8+��M�{QD�c�e��7f��TD�0x�I��:e�^�|���)���������vQ��J(l�n��8����}Y\�	�������޾ ����o��"��)��Tʯ��q�������Pǖ3H^��wy� ,����w؀�K\C�c��u]4��㪆M.2M�~GF��B+�ލÛ��=o��`l�PcPH���%t�X���FW�/�J$���q��u��A�KPP��% q���U���.���_�B�F7�,0'�C���&z�c����JNx��ӛG�&�2���s���g��I��&�~�DQ�ɶ"��P�I�� �X��闩�N�Y��R{ŀ�Y��Z|n	�,�M�Zl�� ���r$��}܇@;�p��_V��Ь�G�_������>y��gV���ɚ�v0�Fw6�|h��t"��m�#�nBpc�K�������q���Ǽ>P�_c���e�����QV�,�&�r�7.�����?�Z�8S���#���w׵��V.0p����<.I����;�>��g�U�j2H:�B<�pR����X|�sW��}���jQ���9wn��h�̋	���'�z����g�oǶ��h(���|u ��qx�2]����\ �F�'�/�}�(Lls�H�N\�i�O�6Ot�5<��OF�[N?���p���3d��|�Ff�\����"(�Ox���X-1{�e�y|1���m� ^��1�Q�X�JE�,���8�cé<�Vz�mϼ�FW��o�^�V3�N��AJnZ-����)E͵�a��oR�(l@�׽�*4�+Mb�Q��y�o�S/�2��஋&��;������0}�DL���*�l�f�V��|�1Z8Q����'u`/���su�K�6۩�0CT55�8���ݩ�V
l����ѣ0�U�Mr(�Mԯ�)�MN�)A�)��9�X轇��K���\�|��Q���G3�L�||����=���
�����1ORG!]S��8S�ە%���I+���09�����,�^](�L�te,���R��n�1�_G7��j1���U�����zA>sp���O�܁���t�-�1�5j@)7�c;J\���:r:��KRr����n��"X�й�|]��_�S��Ej��#hpJ���t��Z4nv�o�Dm��h����a��>A�Ϡq���,�D�3��~}��II��Vm�����;����<��^��d��̿��v��d$՗K6��uɔR�9i=��n��>�1���v�H�8�1,�ڿ�ԝ�0g��X�I�K֛�����$���/���Ҭ\��p��T��E��=�'�P3#	,�3����ߠ{�����P_c!��y�u��x	IZ���wDY�Y��UI�:��?�s�FgZt����u�8�܀�}$*M�7T޴$\x\�,�%H;s�o64�s��.�P�苅����\�R�Ƌ����膖�p��HE�௽W53����w�"pᑁǂmn�0��a���'�A�AF�`Ů�ӌ��Q��y˨~\�J�k�Fv7���\���K� Q�N��9�$�M2�xm/�7� �\3�!bU���S��LT��XDV���JE�$�ds-p��� \I`)d��"�OI��ϑc��̤|����ïRe�k�(�>)��W���T̸�?6b���a16�Z=����H�{�[��E᦭�t�Ά��7�`ʍ;P���_�&�HD����{l����h�r����� z�����ܟ�/�t`��k���`�e��RmEl���� �R�_�jd#�۪�;W���Ea#���p�P��K�j>���H���p�w	)�I��N~0��{�B�_���VZ�5[���,șv$��9d����~J/��L:7��T؃�3�B��w,:�i�Y���à3�@����隢��Ǽl�|b�"&�����H3�'����6�8e�}(���_^��r�$n�_agM�S�g����N���Ĳ�����!~a�pÀ�m�ZR��#��Kz���l�:KKf���=
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf��((�yH������Xd��X��&M���,�Y�h�;�:�ɏg�a���(�F�� 6A|;Ӗ��'���nBq�r&G7�ל4��6��1�]���u}�Qf3��/���5�-ބm�7h����I�r��i�*S��Y^h
���(fʱ>I�y�g�rso�cW�o�/$�A[k;د��c�b��M���E����g��� ��DkgBU5RY�6�1�)	��(T�����r{io�%�ʹ,`=e��C �3{��U�Vs����S�;]D4B[5�v�Y7����:t���Mz� 	$V��~�O}F�CD*�R�~\�3�����I�Ÿ�09����Ñ[��/��
mP��2�Ba&�'S�@���l��	���á��&~�~[��@5�(�N�q����w�P6fT� �"Я|����4�o�R��Y��?��{�%߻�/.�\�X�`
z�U�&7y}K��jQ�z�`�?؞�����XG�#Xla�;%F�8z�;��B.ik����W�!����pb���X���=�#���wf��%����~�cn2�2Ҙ���e"���MBV+�$|/����y��W1���
�,̾tا��\j���Dr�ݙ�L�']��b�����.����]�"se��-���Nx�O��������/ M^:���#냇I���ڧ+�u�JMd��k�i����.��� 4�hK��G|K���W*$��L&7^��v��+@+UP���<��܀3'��1<@B���o|P�K�x�=��5�،�����:�{���>Cq+��U.9cO�zXWj׌��@u|���Z��W���ʳ��g�E��Y+_(��==
���R�"	z�'�Ma���U�H�vNN�(~wZ�"Фf�'D�&�U2��Z�㲷[�U#q�.���o!7�� Ĵrh�]Kj����/&s�A�U����-(��v�����>
�w�!���K�p�[ǲ��5�К��b�	$}���?e�&���԰$��T���x��,Ʌ���I�C�>�4y�d����-���3�=c��>@��o�c��9����-��K䶷��l	�/6.(����?B�0�t�di�$T?A:Ѥ�8x�]?!����pFe��̇���*���r[8 ��!�>����n�!8�P%2B���P�ފ��{�,�Fi �
^�`�k�R�[]s�LR�{=��%k����=�d�q�(��n�x��������Q.��x�׃(1�M�~���!/���+xH�P1�qUI�9"�U���I_Bf�ưEZ�D���s��xWt��$����Jk�ߚ���7�e��R�G���? ?�h�!�}""�?L�r�J
J}�p3����_
Q�	���M2(�@�k��'r�6�n9�{l�1B���:�vy8F��`8�%;�F���0�^�ME����FN7��ؽb s��:^<`@��%i���Һݒ.�Ĝ�T�ȉ���70�r#�OWI�{vYyOe��;���l{�ć}�4|�Q�}�5�5�P�XD� �`c<qmG�I6�gf���1�{O��=9�pg�{��"��H�0ʝE/��g�O�����zbśI��#��QU�B0ʈ��XdYȨ���7P�8�&���a�.�N$�ej*�Ӎ�V� �X�p��k�re u�ݟ3�0�D����W[20�8�r�H>��]pU����^P�[V��iK��&��v�Q�RU��iy�*3���W�v�>��#��d�Kf*�%���y3� ذ�0�;{���
;��������ղ�QC�;Jt�"mr���r-_��t�c⾭�.�#��&~�e<�g>	���Q".ï�� �+�˹=�9'b@�MB�/Ry�g(���O]@g'/ə��������P{�]k��ug�˞㌙�Ѣ���=���y�+,��`������\�):
I:uo1R�F�R��,f���ArE��_㏸仏��]N*�έ^�x�U^�v���Ԓ��MI���B�C��238�|���	�G����<񶦞��4�3����s��è�}l�G���Y��&B\���/�;p�P�b�S��M�bNP$��1ӱ\��d���,fZ���9us��2��o�C�����ƣ!^P���-�u.�G���0�����c��H�]j<��ͧ����-��9G�%/�<Jƣ
{7�+��1|R�Ԇ��K���x� ��'�����c�L��c�&^ )���愹N�A�S�El�vE��RRK�{]���3��U��rc�[��h+�%w����-a�����>H�<x��1w޳���*����K�"��+9,-��,.MU���3�_�)iYuK�Fzl����#��Vh����"C����p*���$�#�z�o�8�.�q#��N�d�+�N��q5���U	�Qh����ʯA�\�~~Xڤ�>[���^�`��ʲ�-��|�,C ��/(S�%����.�o�b�Rߗ�A�ЭŦ`a{2��/h38�ȷM|֊g�������6De�<��ʝ9����rܬS[_(ux�g�2)N�/���I�M�]G�e>RKw��h5-cΚ��PA�[��vW-es"���\�h_��i͠�t�A�y�=>�䜯�|q�Ӛp�d�e�CsY��i�a�G�8�n��PFQ�
|�e��9^�h��̙\�T�C��$!~��9�j{�ήp�a��a�m�ƌ��#�T ����z���gB`Gy��#u�ڕ��+U]�3H���pC5��ez �PJ��j�K�p���,���ߝ8�|@M�#W�Ք���,�����ff�(�s���>��JzevC���V��KM:ƍ��	�&@�d'���:��1:�����;�QkrtX��$�q�|F�G�6 �ʑpk�a��*��ۑ'wr���$��a��:ş_Gߺ���_]��T�#+4t������&G5߿��/N�! O8uG�H�x���u�Ax�:p"��5���l����l����J�����"f �%L�d*5� ���[��*�DR�1ջ%iƠ�d�.%H�
I���./�}��8}�Yuސρ�O'Q�#�3��ՅPސ���45 ��y�K�X�%��{�8�Ǥ�pr�JZ�{��Ƴ5�gEp��4�����ۻ��cM�y�B�)�.6��)���a�#��!N��)�>��A0LqU�/��ݞ~4�x���"R��K�|�"��*u_	��u�cZE�]���թ�?v(1���n��|=� �-)�2k��3�����η�N��ӄz(�F�t�7
	�m�hF��r��ޝ��t고��5�i�n��\�N�����f��Xc,=��x��>�~�w��G6�m"j�OiG�]H�sw�h����9 {��E���fd��R��( �H���	J����Ϊ�%Zb:�h�4C����ue";Oe�ܹʢӘ拕9o��#�P�@�@ݤԧ�6��usr-��a��֪��ҥo�"�ľ������ǎ�rZǃ�ϟ�"Ǎ�?��<��>]K����c[咱����5<g	%![ ���Y�қ�ˠ�Q:��%{jY�=�uX1D�ѝ|T�:����A�eM��Ӕ/��8$��N���_�6/�?Jn�\��(���n��[�� B��ɫڝ�f��{L]5��M���Y�ـ�5��Hy!����۴��1�#:������̋�Yx�8b~S�Rj�����u:s}>P�����Ԛ���f2��*�E�̢�����<5�3e)��#f]������;1]����_�B	�g���W�J�=u[�#bQ���T�OX||'���Y&I�o��|�&��Y���\d�f�����1|{�!���=hk\��*�)���k�ӁK,���W�!Y�)ldPSI��5ZTQ�m�1X*� [&ӞiX��㣫��b7���Ģ�(�������$ɱ�V��e[F�զ�o�<�Y�5��TPЅ,-���y�RO�{�6eʘ7x6�8�%W��<��O��B$r������dƸ��D Qx5-c��S�|n�?����O�ZD.�8]cŏ���7�ڑ�6H��a�,�or~ĥf�ϨW�d���/PdB�]_�O܃*6��ѭ'�W�D^��yV�&e�*⢲9�u�rG�0�S�l:�� �G�|��u���ُ2��g把h�F�c ��zW�3��:��@�Y����O:���-����C�7�f-f��l��d%�V]�T��|RQֱ����>u�q�yCBY^�{��w�`fs(bn�R����6��u����f��!�@��@M I���2�Іq�����~ݽ�Y�A\���go�����#���ɕ������/-J�B� �BԦ~bǳ�	�cNm^qA��e�B��T�̙Y�P��@+*��cg�;(��Yc�le�,�:�����cm��P���0��ڲL��m�7�{�W�Q��}ץ�1�>z�]w�S����R|U���>�)�=�2�̣���iuК�|Ҹ�Q��j�[ؗʙ/0E��8^�pk�tU1��{_6~̪�S*J4_M4�*Z{ԥ���s��4�U��h[�B�K"����r($��pm����R���:����ɠ�P�d��9������)�wۚy!'_�����H���Q�y�s,��C����l��`ي��m����q�ai�{y���T��Y�w���T>z͹I���̙��Vh�Qi�H�G�[�*蟼z�|�'s+��w��M�<�ږ��N}e6}��Ţ�4L�(�G]	S*%��I�O�C~9�]���Kْ�T`�Aߒ�"����Ivܞ�_Į�أ�>@��n\7�_�jߠ��D�~��^a�	��m� -�ni���p�a: �#g��S ,�{&=��/p	X,��k�Jb�8ۓ���#�ߠ�Q�E]2���2��ak��lU_��H�Ur�Y*�8f �*�pt,�^�x�����?�ۿ}&����m-Z��ב�qY�{X�H���l�{����6N�yi�����I�@u�x�o'�����d8���BNE�L�1+,_��4�=kE0�L*9�)���;O"Z�X����.Ns������x�ٽ8�s�u �͆�KU^̲���r��a�F�S�A�����ۋ�0�e��.�'��<B�h��e������
��to���@I�-!���-�\&�	|LF��v�k_ͧ��{q���>ɢ�����:�~��<��H�ˇ�r����ev���)qN�������S�[y���w��\�=i��?@jY�yW��CSa$�a��% �����)����@̳���
�h�%��Bi�s���gad ��5����ಷ0�ۉ�CH??p;čk{!zi����;��/7vepu�0ܡ�5��b'
Y��{TWjX~3�[.l�"�1F�S��
�U��n�����o\�u���h}欺�:�
@�1����ҝU�y;���b�>���ȏ��2">+R���}��عǟ�>dMs�dO��?|�i����+x�\�e�",	h���rw�>&*�/�GҼ��� �c��r/|�4)���h�Z,8G�
<=�t�Ώ�[��}�w&�mQt��Z#�F� $Z�r�r�D`���Cu�-%w�*
%1��uHe�x(r׬z���	3��ە�p���78,t�̎�����fڧ��oɒ�K�����D��Ph��3�;Hw��jy�'���yQM���o��7�k�1ߥ������J9��� T�����0_�B̐��51�S�dFjy5 ��_�'z6#1V�_o������*��.�N�t���U2F��"k�����.�ci�˸}i��x�)��~��������6:���m25���e�-������S���o��@+쌑�s�`l� ��=� _��X�)���C�Os\����ֻ��nP�&|l{��T���?�������#}�NQ���y�e���uڢA)�x{��]� zcԛ�N�Ou�W@LHD���U99a̓3��/)lB4�5�:����;k�$�?�0�[�Tu�<�J!-�x�5��D��d��=�G����fc#�����~.U7�"s�v7T&��g�E�FZ�37嫪���v�V]�!����ߞ�c
A�u�J�&�bbAJ�Р�p2���JS %�6J�2�{����;	 �s'�\�qv)w�B���:���үr@2�<���e�K�O%��Eb.�L*����{����9�Q3,2�ţ�+�͸���<YL4���������z�f
���qm�X�H�0y@��Kd���)xoկXw-�G~���֪��a�xԠ�+ul"�^'��%jH�N�d��E�b���v�Q�=y���M3M7Qs����d�N
X!�_ؔ�W1��1�����z`��JĤ��v�}ڣ^^p�?��׉�y����k6ő����u��������W�t�Dm������a\�Y��qQB3�v%���I,�����ԗ���>:�A�߹ �c}�$sW��8޳������[����fk�7��v�{l؊��WR��"�U9�|�ТB]���4���Tj_�4�#����J����L��Ϡ��Wj�m���&�{��z3� �i��!�Z�8�԰�jG����G��ɘE�x��	����&/�{rxgm�	��|�M�x^fn]-�=����I�̔ߨRO��h��(+��Z�(��GC���q�/�0^V�1eD�$�E3�f���H)��a5�|ce�Ь���}0c�x�F�B���i1~?����8 ڝ`�9�.��6�X.�7�c�Sd|��/!�& �Е�Ⅽ�1-t�cJP(BݵS�{`�6�h,¦���!�����l��s�e�B�Á����n�6���ƅM���b����ܻ��\/g��m5Qg����x\ЃE8��g/4x��;w�[z5�id�yM<�!��R�:�\�j�_��fFm�+Z|�gC)۾�Ȏ\�"@�M8�RI��w���`�^�c��xlw�_V]+��ɝ���)�Qb�	�cлhm��>��ꘑ���2둴��7��ּ�M��h�b���&?�Y�s�HP�һ�������7ҋ:�O8�8�Dg>o����z Jt�O,H��亚~����� ~���LNM��z�51��VX�yR+7�v_:��)�O�F𜻇��[b8jM	����(�ξ8�0F}�n�9��Ą��j&���3�ܐt�oL�",J�h�[8T��`�Ϸ�){�&��.s,�q��(!��n�k����ㄈ� �up�n��ԏ7�ώn�۔�֭�F�e�����6�ewO�CV	M��2c I�{��-{'K�1]�B$C'Щ ��?�C���a�LS��9�w�F����`�ɥ��X��E�{�a�}����s�wy���DV��쾶5-�1ț8o�������g1h����f�p �)�B"�J�L���}��_,uxY1i|�-x����'īÉd�7N������#��Q��i?գc0d }��[]]���zy�B_Lڜ,#�yǐ6���G�u����8����;�.%�?Q�>�-ږ۶����"���H���Yf"V��ɟBwgV�л%��;��$]��2���He�U���hzBAx�Q�U�pZ��b���`�vZ��{�Kd�֕5�Kܨ�D����P���&OMZ(�M�׉GJ�бщ�'	�t�=�S!.]�'�h��� �ClU�壼E;xׁD�0f�s���2��vx�BI>���ћ|�O^�m���^��L��k�����FG�J'ˬN��I.�b�x�ڈT�����x߇�#s"n��٧���u�I�
�]�n���>�ߣ�r��ߞ�:���0F�����%����s�>� { �~/jD��(2��DF�y/���sx$	�C�5}�ع�R�@L��$��i�^r����������=�q�Tٍ�ߨY��p�k�M�N��&Y�{��m#�I �RAH
Xм	zc ;�%sQ�o%�˘"G�}��6a�U0���c�G�+ O8�\aٖ�nO�`�Z
.R�Ɩ���j(r�ҥjB�����=濚�����I�..�8(��#�A}�0�`���u ���<h#��b�>�ˬ����E��71�:��9['�ߒ��͹�B����
���jbFo�/�ZE�������|g�<>U��cd�I��̝��V�֖�כk��8��*���S�ꋀ�>�*21="���mF�b�E�]�!\��u�OtS�+��]����Qp	��1o�%���T���V����}�z��8�Mk]Y��9�]˻���J��6.�
3�
�/1��ik��6n�7<W���D��|N� �����Dp��r�,	�Q��7�*붔]��ͪ���RJ����.�Җ1��~�/4��`X�<�yw�s�R�T�m)�h��+��r�s3�"}׵���!��ꪜ� ��{C��KX�r!�IjQD��o�w2�����$��,X�U��ds`�}=�S6N��a^�x�.����-��5����<��O�%"�b�ȅvG&�z�I�æ�PH��n{o-��œ y��M��0�	p��PEJ�Xى���:�K�`O�'%��;5[�U������+	g��@�B�(9�HM���JG��^.�ׯc`tY�6�tQ��̙��s��џ J��LoPW�\G:QV��f�p$�����h%�j�C�Mu��"�I1����&[��{�./�LC�Y�;�U�f��Y�7��A��w��^k��/R�Jm��v��H�� ;8�iz�����[u�\?5��.�3��C�ת��	@���(�\L�C�Z��<r�c�!0Q;�z�@�r,/�8���ݹx�
���"/[�,7}�GZ�Z��d��Y�����n�9�U��@��.5���yGۻK���ݢ}�Lh\��O���^�43){;뚔-�=�YfD���g�I(�����������4�жo���)W��Ⱥ�����J��0[�)�K�9�Q�z>�.	�)_q+�G����q��[�%(�[;�T���q
J���nZ4z�Qu��!~^�w�"�%
ȸ�x����F��!�r�@tA"F���Z�20����s�lj0���lJu1��i�ӎ�K�qŎ�%ڷ
h�kE����T
�ѷ�����7f�R��NXQ���(��9 ��h�BC
EGv��&��mku�`H[jr����Maf�����,#��J%�-��Q�H�$T�pl:��υ�0���#O����:d̤�y!B�	� _��x���7g0��Ս�,׉`jN#��r�� cY��YpA�-�g癯m�Ҽ/��+{K��9ַf	7����ӯ}i7��8ˋ:�uJ��}�j܎�	���H䀰�-P?0T��  gr����t�{zH����ӳ�ll��ɉ�<0U���D�f���Q�dڇ�GH����ı�.�ͻW�(2�OH�V�UW�ʡ����7^�Kh�rk�_M�M�d]���`m����0M�h})nr��"���i��\݉�;�$AD">rƁ#�Zuuf �Y�@Aifq�G峈v�C�i�;����������ܳ�A���<~{�MKր(� y5yÆ.����*�
3���\���M��H���"Od�$�Hpx[��_�U����(�96��ᡙ�4�|6*�Yw�^�cRφm	l�j���5�hm$�^��*I
��aլ��U#���|'���1��:�3����k��6�S�����\�%�m��q�?G����l���U1E��R�ֈ�B�Q��Ī��h��xeze;3ۤ�B��6��x�<ƍ������;*|�G�?8@e*�5�\4f�����zt���i��(z��A�0���o����ω�1�,,l�����/I����lX�Y������r'E?��O��%�~��McW�\P�[H�
z1�̎[�����y��oOX�n�j�
��˪�3,�o�Zׅ(5�ev�a4$eMƴ���3��Qˉr菥̶�%�PU����A��iC�����m�)>k�*uHw�Գ%�l�b�+,���g�Y��r\����XI�A�q�f����@�v��`�>�G387�����Q���+N�=	7�}}�1�9d)!�v"�������?6����h�>�z�	�N�0L���wy��X\*��Sm����-m6@���-�`2���܂Z�sI�e��>��r��I��a�Qcr�7j�$�l����î�{9jL�Y���fT3��G���?��=2�P��u���(���*M�������fz=���f��%����e���c��.#�����$��~�\�����wr�O�uC��3_��`g�7�+����\)r;�8H1\tj�Y:�v���ؼi`� ��M]S�v���_]��mZ�4��^��2�R�cI��"J�]�tޡ��]���^�y�fUm(f�� ����=g��O�?O1���^!*���*���9�K!��t�#���F����Ѥ�!;��6�4�lc�MW���vb*�f:�F��+#��!ŝx�>�r4��m�~��6&I� ��陻�_��ޅ���i���xѲ�P.��9��������*��0IK"������D(�H��{��d(K��v3vA�o���c6|����l<��Lx�]�#�|F��q8��-"OQʡ�~�=�IB�ϳ�u@i�w��0xW� MM�Й7L��z�m�6��wRC��	W�O:�L�VP2�Ѡ9}(̆)m��(���]	i37�ʟ�}��:�A��\�4L9�Ⱦ���1Ѳ&)��Rk�ED.q���������њ]3N)�Ɗ:����j�͗���ӏ@�ѽڰJ �9��U=`-��D��<1�U]BW]\R �b$o�fEn	:��֘�n����l�":=0|�Um.��a�z�5фj}"@+�#���P�����2�1�f����aә9��v��,������2js���zaf����g>�Ί�sྚ�w���� �hHc�\`IP�ʼ�9r��U���"{^�v�î"^�`�9�-����A�.��j��	�_���C�����y�1 b�Ƙ�RC~(_8^g�z�Q��|���|���r�m"}�+�r�9es�*)6:*yp:���|'
y^9��$��Kԩ�6���]Jw�ѧ�.<�ٌ�ڔ!F�ϩ)���<�ɀO�n�V���ҕ�T����D�"��ǁeZ�>a���c�댁�����a���a�PJ�ƍi�Ȁ�68x�%�|s���	�=֝�A6�0�V�<I�3����r�<A�ٶrV�۽O_����N�s�8$1���3+L�#��1��qC�i����>�ޗ�+�׫'�L�q���5-.ញ��;�o7���.w��|�W0
-I|a�������r0S�R�(��셉�)�*̳��m텤�(���*L��uˋ��!qs�J�6�x�S�5@A<\��q{�`�Ӱ�	E����za� �È���>57�'�� ?����2O
�4�{�|w�|`3L��R:��BG��$�l��H�!�s �nb����FH�ܥ'���U�7��NDUfA��8�J�n��%��	<��δ�z+b����1sD@�"���
0F��!wU���:��}R���/��1���D@�@|�Э�:7	��(���<nn8�W��j�lq�w��[�aO���8��9���Sכ-�=��9�1Q�a�0����:m�Z�ΰ���ˢ�f"����.�x)͂�đ�nf�����}���G�ghb�IF	�y��u?@U��=����\v�^b���0��B8r��u�����N/���X��X���<b.���\���"�,껞�B�6��,Q"��U !�SjfK��\)�ٟ��D�]&���<�1����&1w���7�VR�9#�JUN�w��W�~�3�|R���n��v��TDVO�F����l�hA@���F'%��<�K�?���ʅ)"���yb_���������9!5�������l-�)�T<�������Fl`�@3��W�ܲ��1�DhB6����D���U5�m��飖Y�����[G{��ȻN�r59� ��{[jS搵]�}��L�0�<5��M:�?G�O$K�����N�d�Vj�������3�7t�;� �v��t�8������=�/�s6�qM	�im�Y��@z��=��1ڞ=��XD|�h��.�?�k�0`�ޚ���,B�uPx�=�߂3��1��v�
n5�C i������Qz��ʀ�����HoK VX<E������q�ٴ�%�/��Z����xx���b�xw����I���Y8'w���'O��A�~�,�^"ʓ}/ܜ^�.ۛ��$or�wRV��bJ9%�{`�a�V���[���Bo ���)�Q�*��%���ta��K���FV(�̣�S���D��33ڗ���q������t���#^T�b$]	.����L�F�̕��q��K1�1��S��)����羈reHP�2fS���z��#!a�E���*�o[S6�Q�(�l
j����m1>
�9�~�&U��ß�Բ����u�/Q��o
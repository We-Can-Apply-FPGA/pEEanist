��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�t�!9/�f�=b�:O����}q#�����ʎpH\Ju���#y9?� �y}��8�6<b�5-�l���Y)|A8��'��|sx�����g� �
�N� ٺ�R���L��0��eHXׅE�M��7��o�hMj|O{�	���{{C�J���L˂8D'�Ʌ����%t��z?k�.�l�]�'�'^���_ч��w�(���[g�+���V��6)�gc*�^�`<]w���M���7!���rZF�^U�"f��ď�
d� �l���V
�uS�;���n6�h �S����P�}3{$�=��}�������:��KX�23(��ӎdMm:.JN�����|��G���p��3<6����*c�M.��<�e�If0+�1;X�Ǹ�:oA�?=��F�fd
��ȁ���R駌 �t M�x� ��Y9`�k�ñ��{�<'�%��D��*��۠&�@@�2&>)�)�P��jG}�Ğ�ƛ?G�[����)�`��2�I$���K��OI
dU3�[\��B���e�9�n�r^M]/*��UBNn�	���衠��>C<!w"f��������S����6YѤ�[���g�O,c�{����0e"&7��D�+s0p�#*�k�=�U�p��l� ��ni������R��ŹU� 1�\#u��%��5g����j��J!�6�8a:�R�D�����M����BS���IavB��O'�F�i^�ன�8�d~��V��ZT:��*0w�mD���Q�G�ѬX�mU~+u'���iI���;���]��'���t�)t/���;���jAiؔ��]s��o����X�(����t!��|��D*Q)^���\,��*E���I:zk�k�M�D~�S#ˉ�г�Ӆ8WS앆�4iLc\0�F>�t�F���+��|N �.�u�c���zՌǘ�*+=�[��k�w��P�w˚*��U�`�W�u�7��<`�Bߎ�?�|�k�W69=��*�*�FA���KH��s�h��&.i{Qn�\wIM�79H�=;T��vB;]�C���a��}p�x7U_7M����$�=��IQl���HA�F�K��=�;���[���Ã�i@m�؂�Z�os��'�;���T�5�����a_�]�.��WmzD���c���j����|�M���Kr}�����t���թ���:�B7�F����Wf�<�Mr,��	H���i��<�_Tӈ3�q.��K����^��sMG�FO��KD��d�,1��lu�4DwS7Rl���+YIQ��+ �&z�B�?~����	��v���,s�j�pU^��ě_��_TG��?i*��]�h���_����>Xgi���\2���^��Z4��* �x�+}"�E^A�q���1�r���G��5 ED�c+_e�h��L�4!����������v?�p�R�/]������١?�^�R�t���jĔ2���AnʂG�c�c#cTvf��=+�Ҋ�^���B2�������(F��������a|?=y"��i��&�� ܂�w
0�b�d�e���'n�F폾R�$,�����TUy�m��:�D���SF���Zg\Ij�����N��a�����L��q�(���k�r��@�f�,��p��[�I��gڍ��m��
�����Ï����ɐ��elP}��y�޿W|����'V_5�chv���ϒ��C7R�{x�����	��T����L�e_���\�Ns��R=?OGcT޿�,����<�uY[H��>@%q���5�n龙�j��{�l�5*���ҥn���6YK��\��-�����"�n%�f�:*�>@zPE�@k�f ��HI�B�<�_� �������y@5�F���)W��W�M2 ݂��..7��ʀt�R���os��r5��Z�{�����9�S�,�1���mA��o�F���.�shڣ0�f���gj����X��g��厨��4��5g2s�3�tp�e�DL��J�bN�pmP�?��\�p|kc���T�~q�Z��)�!��z��S�몑l��+�V���,���!T�D���[]ä�ʛw0�<Q�$���+�a!������=��~��u��a����B���A����n�q�JU��g/��~��P���
[�m��IɊar�K�Uf���eH�ӳ^rw�D$���"m�25�?ɧ9��j�Ű��?y�@�<���Ȋ�с��/�I���l�i�L{�n�F�XdWQ8�u_wz�f8Z�'�bH���dg.��(�	u�u��!���O�"|!&�[~��lO�.A�}��0R��,iLÏ�� 8YAg��Y���D㜦�kU���h��Z����3�ẃ�.���RٗJN�e_�W����ݿ����Pȓ=�	Y�.�֘"Ւ��}T����d�k�Q�yK�r��3���/��?�h���F>�ɧ��)�e ��Y/{$m�I9���F���=������Ը�>^Ʀ�v�$�&H�R�*��,c��~VHQ<�eZ{;{�MU�:�D~_�_�s.:$����}�r8��f�˼y���A��M����=�z6�"~[���M��k��L�iy�x?�!�5��<QQ7hlW����c+�Vb�0֔�+'[����@�q{ �ue���̥dr��j���� ��/R�ϠdiJl�&�v��oF����<Y�e3�Οe8殮����I>�#���M�Ȅʖ���^�:�+�2�5�����G�Jv���>��T�u�9�Y��Qg&yA�aN��D�5�I���|�y�krvn��{�-�	X������TS���٘e�u{�cHG����0l<��Z��j�C���0ь���
'F��{Wt�Ș�Pb�y�l��P	?_�sW�՛*��G�xWi7$w�:$6��gr1y�3&�ڄ<��s����Qϼ6�����j!%�p��E���PE�e����C������U�r��k�C5��L�b�A�\���?Md��
Nm�t�/��rB?*r{��>���.��
�l�9�*���/;��<O2��-.f{���)@��枂��o׸��%�<��%�"M���u/b俀���op��S��!g�ى%#
ջ�A.�"�)#�<2*�b��#v���4c�MD~~�-�'��$G���v�j�%�'��9K}e����w�^��I)˷/�����D�=�E���g@��!��f��b;�:�d��kHu�ͥ��
f2���T��<��!�S�kb��V@�%l} A���L�L�Xn�g�6��� ���䞸ŞN��7��O\MK�掊*5�$���i�����-��Ġ��8I�PǨ�o�,&��Fq�,�)�s�3��}|���9]�Z��V��Q�~��\�R��������f��Z��2*�ykꚚ�kE�Ӹ����@�)�Ȥ?r�{�,�I�s�L�m<֖��|�&U�ʆ����<�����C�9TB�^ݯ�DNq�x���J4O;��U��8����&���;}ۚ�%������*�3迋_8�Pf(v�N	&�I��d���o� z�q��b��P��M���!�@J����E�S� Kwݔ��]a�UbU9ؗ�jf�jH��ͻ�h����x�}�MT6P�\g���2�T��Q�D<���U�~���]������ %����]��}�����Jޏ��j<��+��~=�u�Q,��*w���pQC��h�PGBs��'����6KU�C^�g��(V7�m����)uxP�[��F'D�N�p��u�9T�9=�ř�e�q7�!Ө�. ��oU�9��'t� E� *&�(;�n-fE-�i�!��՚�<���j�r<O֯���a��+ox���-�:��c��AwKV�%H����r<��W�]"!�	㤙\����,�ƍ)���N�lW��[O[����>.Ĺ�ˏ�����������4�A�┷�t�:8l��gG�$��Sj�?���k�@�1�X`��%��	��ꔞ�7zW0 �c��!>x�`7,`(ٞ ��DB��}�kHP��m6���A9�V�9�$d+����5:��hUHĺ��A_��W�YQoG0z?0���fG���ΪCs����R�h��u7�Mk�)��3��}2�Y���e�^5�4�%ZŽ�]��N�a�Q�'��.(��3�	T���:�,-E�]%����9��,�OX���+pT�������3�b'j�p
�>�hV��Ũ%a���M�fa�?Fy��B�B�N��L.(�οm\�.n���h����%>)l;��Wd�dT�W$6��@��r�2[gw
�{�e��tkf�!^��� �>;�>p^Z�%ϝN��5�f�F��5l�)uWEO5�I��ݹO�)�c-��B}Xr���Abj,�Z^�x��+�`4�j��l\ ��Fx�u��� ΁�ę����Xfp'>&#�C
�UX~��<�v�iSp����'�{f���t�'��R�Qq"	��L��!R�v���~e�J���9w1���M �/1L#���r�+)y�e����"uۏ�/V���{���@}��]���=�:5t��C�m_yĬR��;_7ؑ1���5Ss/հ� ���2y!TƬT�(I�(��x�+T����͋��bv���3G�h�q�(U�nI�M�w�;��%��`�.����������͡�ݘG[�iT��~��}�џZ
s�J&�6��5���ݔy2�GP�UȾ�Ϭ/���9�l.$����ω��d��7GP�lT��[Cp�Ne�-lR�����V�(5�� �[:��$!I -Nֱ�알�����v4���&�w��hOT)z�M���Oa�m�K�����ǣ�V�q����Ē�Y�XD8dLo ��vBV��K�Dwo섃Ӳ�5���!���gG� [����
��m�H?{C?J��ϖ F4S9��-M[����An��^e��C�j	�2y��6�dm�2G �	��$4�	l�VeAh�_�=r�҄���<T��$��q<����:�	���I�~�CȒ0��ZM	»���2g�R��=�����=�~2ew�9o�c��|)���t%��w�I+�=DT�C��=k�D�x@o�k��/�������>{�z�g{}ōJ6�
qn�d�m+�؂��C��t_
'�=KC�H������� �'���ּb�1(�hE��JA�:3����54[��}�S�߶�/M8�,*�0.��:�]�[��*�ѝх�Eۭ�bI�nGߊ�y$PC�I��맠+@}����\	`VZ�
�?�|&^�����/��IR��Ǻo�Gx�7ò�n�`���OZ��Cצ��z�@S��5�b���%��Y�p�hJ;�|��zQ<w�#����o3����k1���f��2<-�FP*B_�
uP�/#���9*�jO��\dB�هp��1����C�W�rU)�9܏Å�׽Y2g=C��)��^gV��Z���I]���/�,p�#e �E�P�ci���X�kGC�Q�5N�xPl>�2��T�S4&c;K��.�"vb9��.����=@ U{7�}t����s�ԋ~vn�g�����A��w7t�/�͠�»4�ZPb���L	+��~IT�ŶK%�¼���PcOIg&�$���c}�Fz�S���.����);�D�ڬ�R�(뚯����=�� ��b��S������v��=�f(B>���S7����F��:7�1w>ba&�[�E��5��h�����/<H�9��E�S�)�G�����˅
X㷧������t\�A�/��]�)��5��:?a��k�Z<*�_u�!�0�_f������ָ5'�(v�QJ& m�E��r��$��P�K��f��M�rS+��ɡH첸��0�>���{F����O=�;xc�'!�A� ���x�u�o�S�}�9�q�^��P��И�Nt>��J�r�����W���K��+w��Ӄ�ڙC�X��R�"�>�a^�e�Y�X{�(�~��L�_G���n��Ih��!ҷ^�,C���@}p�&����uGU�Ζ-T�K�-�i�f4��F9��"�D�����L��yߠ>�q��� D������;�e��:,n[����T���K{4��|-�Ұz{�\��b*����j�	7�C���M#2v���G�Y k�V�Z�O�:�]u'�ڶ�/I�&|G;��%�%�s+Ix�0���䈾$+>
BN��Q���b�	� ��
��@�VBE��}����6E���.��E�zNF����%��\�
j�
��� �~'���C�-5(�y��,Ho�qM	k���{,?�g����qJ����`X4uV�$��bw��i�����N���.'M��Q�i,N�rf�x�3E�tÚ�����ܯ��h�/�C�
�q�s3)5�4���zQ�4�&i���X+_����Q��[����v�J
j'9�7�CF�5�Ep^���1j-�S�L����w̪8��Ƙg�s9�Д��3�˲Q���f�%^sR"�PD=_�0�<��;��~�#����f/8�"�?�R6�:W�T~�+b{��F���_�(�����8w[d�k����O�Z�x��\�ɠ���c��0%��Mr�����j���b\&���L���u��3��R"�3�v>/ǌQzb��8����]ZR����ڄ��ů���i�n'���E }+��=)T���΢fx�V-KV��d��'��2q6�[�_��b�9�0�J-,r�|8F��(�0������io\=��e�J˸JƓT�����'�V9�B����SQ������!�BG����֘T ��[Hqv( �<(v��Y��.���8.d��YlX�D�� ����q!V4��#��;d��T&w�'$|�E=���:��l�q�/?8n8e�MQOU��H�����/��bC����B&���薸�G��t�--����6v�������-_�{p����Ɍw��V������E=�0 )��3��=�r�=!�����U�t܅r��~�z��C�=?���w�����U��ChlcR`i�a������T���I�����(�Ҹ�)�D�8���1����Au+�l*;����^�[�;��&Pz���X�'z��p�8�xǷ����.l)�M���rI��l}�N4��ջ5=!$��,OG�<�������`��#�l�[�n?�?�Q�3�HH|�S[]c�������s��~��9����@�w��Q�G��,��Y��79b��mDc�'Ɯ���ܶ7�e�]��/�~�Jco�e+��&�t��{��k����� ^J�� +��(]��}*��_�T�i�E��S�'�3uyu�L���u�VA�����c��NݥO��V���>��	��/!�$N�X�mbI���``��<h����V����@�W�J��#oӂ�����;@�D�
�*W�u�'<�V��A�]��a�����H�ܚsRf�����2_�7�;�&@Z�[:0cf�ŴX��:\�&m�u�g�@%c̿/��P�w�sg,�fԼ"m�D�蚁apONs,k<h�J"������Wk8.շw��B�$���S�A)�C�BJdԔd�+1 9�mUUZ&1�8������C'��,��|�&�> şm43j�V���ȟ�Xm���w/>Z�u ����uv󰲄�����N����q��9�% n1�^fxn����wI�� ����>Jܩ��H���?_����'Ӂ����.o��f@!�Fo��`MT�cnS��c��"�B�(�W3r��`Lȑ["��\�x��/5�:���ǡ .�_$1RS B軿�9T�7Ep��{We�V�: �Ʈ��ӮMe:!6?�h�,�K�Θ��p²�CMb�������=ei��+Ў��oL��J�3���5�l@v��k����v^q�D��mÊ���Ɏ�@$X �pD�d��7��=���[Z�m���_|-^J��dZ��U_�_�p�@�ulc�-Z�k�&���>ʧ�������+<_�p�V:u �U��5�6��9�6L��o�:ϛ0�cX��ː�*����~�ObY��z��\�ݰ
-���e��a<H#^�QwV�uC��3�6�pI�r��.=�0:���@�Ł%�w l�L��Z��՜��a���)���Zmd��~Ց��|:�{6�j(��)g\,�l;DxZ�[G`8�uR��O�`\z�`?�����b|�r�`#����x;>\x�^Z�~�܎Y�)�".A�n#��엂����+a����N�ϒ��^�X�	�e�<�F<=��5��e�,&9��n�P&]qģ�j��mj��d��M����	��� (泊b�Na~H��0ʆ�fa��T�wo���ב���z�D�",l���dؗPj�~F���$��$�*I�]N5j��)��bRSf����>;��B�fB�Q�DANE�+[��=c��N[��i�Z����#W�\�-8;��d��R��$��\ �0�f���Ю�H?f ,�<ܺ_�����vlfr��	+���(��91�&K6�H�F��N���BN�xSJ��+;�vHjB1I��DI��``��vP�kJ��u�QC�.��ZɥaF$b�����k8K	��BtnWUaC�]���s �߽=l�����ܯ���`s(׏r4�]^|`bsE66)�{*���Qb����$����oM+�Ov�稳��R�r�(��/��k"��_�F�Af��C4[*N;��!�Rbְ�$e3��p�g)9���J?�u;QvV�I*cl�J"���Q�i%w����ͽ���6E~�[)��o�������(�%& -eDM��Ϡ��?{��Gم\�+����9��<b�P����D�p�0�ok�K|�x��E�nZVH��B:�쎢9�7�*�tn�W�6�����(N����r8���V�c�������>�8mtT��������Un9�: E�k�b�5��Gw���_@��_���Ơ��z�Xؘb�A_8ɵ�n��G�û����Sd�	��ydO�G��/�C괴�_m��w�x�
��� �v�P	�F�
�8e6�����
��'ģo*����)�=K���mb��j�{��-��s4y`��0�^Ѻ�n�Wr�*�R��J��Kn���T���x�{�M�bn\�l���}{�"�^��g����ϸI���L�ԈC����?��3�S�4����!�F�J����Q��Qc�@h� �0�_���Mm�h6m�fBJ\�fdbZ��y��1����ݐ�	�3�ZG$Sk �E�C8�5W����ў�[O�vP�ϸ��(	[r�f�Q��Ҟ��K�f𥔚� ��X��B��C'�ޒ@��/3���)�ݜ���K,��jW��-��E����Q�����HI't¾5ՊǾn�8�s5a�`���=��y(���4n7Z=�����)wG�D�F>���FހW��3���:�a"B�:�PsTLT��obV�G�`���i��S7����-��Բ �.-j��\Ȫ��8>ĉ]�Y�-
G��e���	��eL��[�G��x�4pї��=�M ��w�qj*���{?�z�w��m�����h�p�q��d̦eJP�g��p"���+2��k�t��7�n��J�����d���F��h��v�@�/�mPlY��	��|hyD	颢�����F��X��J�y��s�@�Ć�7K�~���2*��)L[8"�������H�$T����q�xML�1�m�dY��bz���4�C�>���݃�9*�z|���as��9����,��!�d�iS1���,�ɞ�I�P����h���5�i��a�4-Ks�:̆�:�v�u���w]�V ���$��jh���g[ۀ�A���x�|�F��v�Oo!np��t�Ͷ���ߴ��%�Ak)m�Ev�&ח��,d�(=���P�b�y{z����l�2���*2<�{DYP$�%��Y�z+�M�:���e�ڜ��3Q�X�QC�u�)��<ր�[�_9ȓ����Mn^�R�+�+b��Y����`%����eᤚ��l֩�FH�+2�7�֌�s�҉��$`���A�x�Bơ�!ƅA�>�8%̥v�Jݱx��p�t�=R�����+����8{���tL�.��~o��0&��19�r�75+�UJ�p�9�ܻ~o�+���~�Y�T����������@> �A�E~� ��d;YloN0$� �u��J��`o�B;�(c]P�̪2qY��O���=�> �'�r=\�2�*O�o�O6T�Rw�#͂Ov~ߔ\ r�ÔG�L��F]����3Ô�A�H�
B��c �C�=k�ր9�yq(�"��N�|k�1k��1�?�����z�|��J��m;ۈ�W):T�(��sPJS+`�#)h`ﲺ.��erMWY���M�`�ܡ�L����=s�J�c�N�⮪E�A2"Y��NrnZby�`a`8�)�AxZ��>6\�|j"�@�)�5�X�8n�3��f�ا��?��"���1%s����Z/�Ќ��Q@�<��Jz�ejb�S�7��y~.�l<`�#��e3,�C
y�.��C�(��륦����	�|Kް��K.����Sy�N�ъj�����-���(�9�L���wԷ^sh9�mX����=�pAv�5�b��-Sw�1Ơ����M�<ǝ�6�"��c4yx���ue��K�pK����D���${������||7�D����U@������O��+Q�zo�ղҶ{�<�r� .9��u*��1޴����#�Āq ���ń�i�R�Ѓɍ��ߵ��#��8?�|xȧ�G5T�>�����$�|t�K�g��vig9�M�'���k��s����~g�D6g�W�D+<זg��z�*��^�FX�VQ�=]Mu�?g�l���|�Z�>��V��_���`⇇d��Sip��%'�z��m�{�?�-@��m0�4t.��932�F�V���ׇ23A�es�'%b���I;�j��cD�J��%;I4A֕e�����9D�}J����ڷڿ�<���%���d�����7+?�^PK�3p���!o!���*��sı�&�03�>>Է�/z�Ǹ�����>B8��q� �ã�`�G���L$u8$L�2�-N�.�$K���:�eUv��s��Q%.����u�_�[V�X���} �?�L�n��x㹦@&5�iI񧫹r�]�1;�g|�ww}�h�g�2f�]�S�-t��-��o����
��6�AH3@��=�#�x9�����V7�3T{[�N�k?��ѕ�0��t(��\D�����-�\ug;������4|w��<�$�N���(�q� #t�R�O������:�VJ"X�Xv�*�{	�n@�r줮#ϥ�6D�8I�?�=��:�B�K�qlB~����8��voťӀo��h.����6�0���d���T��7v���z�Q���p�UB-�����,{xe!�M�}I��r��?��*����m3�t �+�^[�y�0�*TLmV�s�%q?Qg�<\��5?��A��O�v��l����h�Q+�0P�a�f�֐�Ҧ�ư���o=�� �_Q���)(X	4�O��~����G��$jc�2����b��ue)ϝ؝�k�Vf]f'[M���2Ky)�'�_)�"�v��d�ȑ׻t4޾�
�l5e���#~�s��t ����r`���2^E!�1����p��Ʌ��KC�М�Rw⧲ꄙSHQߴ��:M��Y�O��Q&����5�󈒪�Cu�H)�Zf#��R��q�� �Jq�;���_�S~��S�>�{f:��9+!8EHJ�(��zO`P�t+��'�{��	`9+�dN t%b�}�&r����jJEa��r�;j� �&V�K�@'3�!֡߀28��"�aG�j���p"(#�TE�F��c��-XΒ�q��ޑϾE"2�邴�VH #�L��}o�xvQ�Ko�W>�k|B��.���c�.5�ӻ�G�X��U;jq�U�i�\g�h�+~�Ӏ��b��o+�>���t��T�������)����L��0̑A��s&��I�����[8d-E���@��Eq����Z�Ҿ,/d�<���ߘ��ve�����n��Fu(�i����"�3��N# ~�����XY;��ջY����@&���C�I6�8���+�7i]o[���(�#�%z�.�;�Oi�y��UܷGw\F��_�f��)�u��AH��,/naD�@1Yl��}�b˰���O�{Y�}W75�:I����~W>r�
S�U�Ϻ4z�G�!̿���+Ood�k����֤Z���T=���81 ��(�E4$���G�,�Ln��`�X+�S�Z�:��������D��N?	$�dB����Koz�q�F�Ql��cL���@yW#�Kt4_"�U�B���<�<`���izdԇ�/��cE��+a�3?a�;��"�d#�N=����l�K��Gl���fZVe�yRH�R�aSAՍ��2+gP+e3���Z�F�<��xwO�@�`�~�!px�x����Q���D��0Y���&�ʖ�t���u$��j�[�>�G(��"~�YB	l�4\2�䳭�9�c��ri�Q5,>JL����$Zo����u�3"��07�i�?��J�r����p���5��BU�ʟ�H`0
͆�=
���@�U��7w�	���P�^��-��R���c���9���U�ݲ����n��!}�%���{e�Ĝ����zs鳾���'E�R5����$�~��\�Ծ�ĩ���X���W����-���O�T�±�nS�������ig���rB}A��?B,���}!aT�#{����Jx�'�wS<e�jL��� <<�m�u�9΢�/IS��?�JT�X:�(X��@�E- f�f�o����q������$M��H��%�BҎ�E�ۤWc��ZDVq(h-����F u��S�M���w�d���RQ<	5H|a�k��ΖQԻ�=���r�?�����O��8n�kr�����-2�ס���]G�`�Auv��t0�d�	����^G�P?���SX��:SW�{L����U�W��g%H���t$z!W�숻H�p�29�V�}1�	���;Hۥ&��X�g@��E�b2R��28���A���������ΰ�a�i!3��fܓ�Z0�~$�~)��;j��u�emCLv�^A����p��N
1�}�s>,1Ԓ��9��r̝��X�r������(HG�p�2����.:A�=���c8%�p�
!����Z6�ƣ�7�Y���|��ם����x�RP��<d)&"b�_4��ю���N�����>nrÌ���_0=��rj�k��@�8�z@E!cRHP�N"`�Ȝ/�r����ρ�qx96sY�T�ф]�wc��lY'����j@]o�v��\�
y�����a,ӭ0��uۿ}��('���a`\B򭼏���v<�#V�N#�c�X��c���_;b�=O��y�� �ў���o�L%�"�ݡ��P��>KU��yuZSUԹ�
�0�q���,%�4�o�@1uL!�
�О�|�0�����A�����np�^bG0G�y�QC(�鋀6�[���j˟�7�<�ėB�|����E6Ϩ��4riqX�!�
�>P��&���	��ҦA&�:<��{�+ȅ`�%�Yq�8���5tEFT�R࠳�,x�㛔91Qjn�H&��u���\L�:k(b��jD�����x���
f$/�����¨���'&��پ���^�Z�N�LyK�j�n]����8cE �u�Z�}~�S寘�7��z�
1�,�&��p�d�@,q�����2ا�� ��-��,T[��v��!@*=\�P��+]��}^?����<�7D�q���A`�y�E�m���B����r[0E0N[�\�ݓފR���6�e%�a��� ����Vh����<�V���,;F�>�ݣ��E��is$����S��ۺ��)	ӕ� � ��`A��j�H�����&�b�YkH����GK��/NdKj�J��`�hi⦌r�}o��&wך�Y�a�
�W��^Vv󮟇����/�ҷ���UT�`��{8,t�D�����k�6S��S��%�l e8�����C�_[O4�*>ޞVv�~��];nn����(���ݓ�(�V+�j1�:��[Ix��^�����l�HCY��#*����U��W�y4 MmK��4s����c������K2ޮ�c�x~�l����}?����׳��¬�h�Sf�5װ�4q�IZ� Qs�ԻY��gM!�qL=�_���f!W�p�-�Nq`�����;��"�n���m��)ڴ=d�K�5�2����d,��Ԯ߾�J�u B"D�����M�s�kXi�X����4��/�d(7�GhM4���-��6�v�~DI��`9�XK_�[	8��DJ.��vl�h@a�la�#�:��ab&:��ˆ�����"3'ۼ1���� � T�=0`�J�����?���5y�ڎy���� �e����TjYخ��7J-�z"^�/�D�p�N��sM�JӋ�pJ2�S����fg�+��:�	B3��Y�=�Js� F��Wm�zv����P���DC���j{�Y1*)��]�"S��%�ܜ��Y/�֩{x	���iL�Ug�#
��/��8Z�L	��Y�@m�@O=�&�c��q���׶�!��b_�@=a��a��A�G:�w�DY�4tG�~��TY +:�q���=∛D�[��SM���q�>ٱ)� 4.Y4A
,��o�}��F����w�N�����0�e+N5]l|���=�o�v3oTsg�;���
�����b����m�-�s��@2\����gU;�N�p��
�F�#y$�[å��jY.�Th���"rn,)]p�'˰���<�r��g%����h$`T�"��z��i�����v ���(Ou;�Y
�\f;I���=�H/̈��� )��֨�j&��>9�kWi��0C/Eی��pvC��2�L�&���h�^��	裠U�])f�P�U�;#�+|"Qa��m�Z�6Y�&�j�pn�t}�L,'��؈�g�2��ey��a��9�繣;�7n6 f�M7Y�D� 4�R�l	*ױˋ�$3�G����-i$��ⷩ�rŪ�jk�\�����̎�+� ��q��� ��{�`��h�oDN�`�|�)ص���GҤq7�23���N�6Bk�*�C��qq[�*2�V����}����b@���5|�A\G|���"�E1���̸0@��V�PP'�?�_��/w�ݑ�`4��Bg�TE�P�-�:�`y!��[��X:�=p�$�[���~(���)y�]���/1���k�@o6���Iy��8*	.��t��;Д����_�≦V&Ô�4��y��(.%����Z}��w����	���&�?^~x�~O�G3m���t��������r����e�^���۠YPg�k�7���D
mތ�s��^&K�s*Z�C��ͩ���͞f�y:�������h�Ŭe��݁�L��AZ���{��r��z|��o�Z+r��Wm�Cdt�ᥩ��iHK�d��ۭ*,�W���$�I�q��>�s��r��Rݦ7᛬-�Ap�;���Q{��~@�+�jyzz��)������K�����xa�t ��<�=���g���@�7sк��&{�;��A1�i��Q�tG-����7��:�F�����gZ����L� �a�m*��_�oY7{��v"*W��<����˽���C��t,�T:yUK�z}�X�X�;�����n5͢:���ς5����L��l[L|f��\������*\[[ߨ�V�~�<��6�3��L�I�ղ��=H&KL�Ȧ���f��&�Y��x!��-�B�T/� ����]�d�F�s�Y;3��C@j<�d��s��<�P�y����z�"x�1Ox�A.a���a?%t�%���G��R6�ߏ�����rAȗtx��<�?�^�����l6���P��k���^0��}�2����Z���pR�Qx����CE_�M��.���m�X3���bW�ޝ�^SR�3���>��w^\�rh�
0a�U��K��r=�_&��7T<���87������.^BU�SP.�5 �B���a���f��Ê�!_*j\��Y��N�,�S��]���\���j���pco��D��9��	_1~�_��g
�Z��-A���N�V�!��d�*P�ƨ�4Ҷ.� ������6�[:5\d�7CJT�g�Ϩ|nMe9g��"䩔��*���N�?昚^������$qJз|�YT�̀��T_Qe���Mt�6��U.�m^�I�9b��CVc�|��:'d����̥�Nb"�.`�+7�w1�C���ړ��bă[%r,j����Vz�Zx���}����=��r޴��OnH��CN\�V�O����ݸ�0�p�=�Y��V���Q�t��F·��N(�-��v��(tg!]��zwKT��>�ZihΎd�.'�������Z�,�������r%�R�e��'���+r��f^z P�&�)Č�^ğ�4�&pʞ�F�h��V�:�뙁:���2UL�l�8�[]?�g#�"�j�Z�3*���8ֻ�8�}��3�
6���i(��x1i��-��߲e�k�8I�Kj��������~����b{�k�v�;�ZlL��?�׬r�/j�����,>9X�X��\�M�<���"T���|��s���i>����u�燫PzC.�^C�h����@
8����]��>���  j��.Fn(��:������)4لY�:��Xn\�n�<�-�9�?̥oM�҆�֝�m6K*}}��1��&��Q9�%�.��{tSb�U5�Hj�"Q{/׆��|hhS2�[��:+��ÛV�G�����D}x� �Z{����[�e���L�"��� Q��!���֢4$"B7��-6�=�98�
�����_���n�>����M��%�o}�������oJ�hA�7�I}�"aɭp�)�ڭ�����G��M��@�܇�T��.����kt���ai���;�j�al1A#�e�\.Β�Q5�FEH��3=ݧ�^S0��
�t�GCf�A�S��9�H@
c�	���4���"VIĲM��)�� s,6H'C��$	h��F�H��Q'��o坿W�g`�t������O���1^I%�g��&)�a�k8oh�Db��m����96<4|M|f��:�L`����k�ZV��$@����ڳ���>�g7qsYr[���Ƹ_::u��E:��+���T��ƣ�x
?�#����RA��
���>��+ (z��1���{��,�x�Ԗi��R�s(��!|�-�dXdExR���{�����t֏ ?G�0B��e�B��G� ݴ᧾tw�X�l��O/���.���ڏ�x;�Ttj�w�擑l1O�܃n�W��`I�T>���K���Ia)���0N���x7��N=���2c �@�f��U�9�PԽ~h�.���ܷ1+�6�Kjd����͙�Vf �رz��;�%�;�sS�c87������'�˙��R��<ҟ�d"� ����F�\����bv�u�s���T-9<9tz79��k#\T�#�9�DF�{��2s�b��)������qʹ��A	M��Z��ަCa|R`�k�b��8hF?�,ߗ���4���ʈ,���fU8�J�N��O!Wa	)U~�:}�In��9e�պ����Փo���&�*��dB�~aK?��{Δ����o��M�^Dj��\�G�#~�_gE��P>�YmV�m��^�ܟ�h͠ uMz�G0�q�|������ߓ� Р��p9������|�tI��@x������6��>)�z���X6TJ��.�)�+7�n���t�r	��\x&�t��k󃵗�chs|������7�+�X��j��|���$��N��8�)���b�8�Q��5�U��(%�Hۀ	����9�8���;ŔN�7}��IWZ/�E�✻�g����p@k�Λ�}؉�o�&w��<_�v?P�D��C��}B<�{Z���t g��2�>m1��Ď��z ��,�l��Kp�8�E�ɺx;�I����A�E1BXZP�d�SJ	�ؽ�!�Γw��P��>[�<�L^rS��8J\�H=�R�s���Ɋb�<)�;�v�[�f4���ΎZ���������x"p��d��F����Yx�Ul�:��h������V$�����A�pU,�S;�c��݂h�������@�1�6w��Q�R��ڊ[��?��{� ���|����7�Kc��4N���}bXi�M>���'�:�5�bS�y�P���J�d�7aƙ�w�%���!�%qc��;X���\��+�{i�-�y���#�����;���G%�+��'f;eK�܌w��~mr���H*t���>6�5�KQ G�Å��%�}��G��_:ki�װY�t9�����
ȯi��K��r#��4!N>`�B��usN�	����Ǳ���/�C�u�'�6���w�*ٖ�u4�����32S�̃Z֥��}{D@�^����l�<aK�m ̴�,�Q���L�8v�S�M����&����*�(�mIcLC������ȵ��㒑y���AϻW���cT�<T��\�m�8�8=�ըHl�V�(]X������cJwg��o[|���<R%� T�u��к�2�W�ݡ��;��f���X����KIg��n�{����� ��uֱ��8#K$�U2@�	0v0���Pt$A�?a��`���� +����-B��\85�@QT$.�c럑^��%q ���w�Q?���^^�ar ��vH%���Vů�9F���V;Jn����4�I��<��i�w�J�笙&�jS��:��9��tr��ʝ����	B!"|5��(�`!L��ۻ��$Q6��>%�z�AIH�s��9<h��k)P�c<CS�$�Ǟ��o�mcNe����~��4�8�?`���ǟ��d�Y�yڤ0X>^It�]������FC������d�@ʳD6НYX&�ƳX�?.���ie֊�"���ǖ]�_����LH40F�u��_G����]�/L��nO�D:M �2M����%I�pUFL׭��#�O`�xW�솻5f���)W1�� �P:Q�hѓ��Gs���!z�o�j�hZl%O��6���å��ؓX������U�p�m������D{�-n��y>*��*;�[*V�jE�br��)Zq1+Sq�����d\�8�V]�1Nlee0y��j}z�e=�)���X�S���h>:�?�iWY!������L�ų�;~�6J�_ۘ9()������yߦ��?4i�m��K8����ҌV�j�ֿoQ�S���X,XG~�p����}D��g�6#Iˤ�}ُ g�/��W�=W�^U��I)തB�����XQ�D���W��ڹыi�	U��0[\�e��*�,؋���9�PH5g-;~v���UiN-吴�d�+	��3þ,�!ˀ��s�)�3�'{�|?�l�(��5��ob�![ �4D�l�*XT5�'�L$��#c�
���pW��8���2�Rz'K�v	�����t�uho�b�U��[��bk��ڏ�>7x�j*���'m��bSz���3Pҵ�������7�%���B���oǞ�]�Od��0sG1�a�����t��wdK�*�����A���-u��7� ��:e��t�~nᤜ߲B�	c�$ۅ��7��Ă��azܷ���?�����U���sx'��SG�f�ɓ������"��u˒��YUz��c͢�p`�B�	5���_qR�[цp|�[��Z�����1&��w�uLZ�S���nV�6[�D��]�J4���&�ߋ)Q�n�mW�2�C���,�c���}�kD�i�=v�Ҩ��aKS�1�5��B��F�0�8��:Ts1��I*y�Q�wؖ�_q�%.D^ms�����_hd��lv4`ҔE�T�B��ćz�~�:Ԙ��z{J�[S���V۟Ms�,qm�e��RJS�ӛ�k��m���Uli��pԵc�3�N%�&3�#����g��UQ;���0=�!���|�_�p�׍:d:ó6>�ӵm�	��@E��!ڴȐ4]>�X��6U�B�����T����s�3"��X�n������'��̴�����)���o+���E�	���/D`�J\�������5�G:�>w�=Ch��s/��B���K1u);(7qkY�MȻ-d��N���x`ԅ�r� �A�ŭ�L4���J�V�@4�V�]�h�VH��*�Q-�!����ԛ���F����[K!��-��P7ې�:F����jy>g�_�����v	'������?%�����ʌ�ݴ_lO=v|�˘2��N��ޱC�	~���~�S��x�1=��X&)������w�~�a���)>3��i��c�g����إ�Z_����/#����ʮ;���1�	�ׇ��7�R	�#_����/S/��	EvG._����Ԭ�#Й�:be��*�������vFQcϪ+�FR!*L4�
���Z�8���B��>�*Q�{B�k������	��]�rD{�Nf]�U$�;��zՇEK0m�� Lyr�$������u����K�O���4U��`k��0�
C'iG���%���=~���������	�� �gI�hAx$�L�W-�{�����mV[���nj� h�Ul�,�K���
�8�X����LD��S�P��de9P�fZ��������$�xl�杒kcJ��߰WF<d��Dc�J�m�p5 S��,@�^ �8f��G<��خ�A�SOM�V�_ɽ]�k��>ܐ��߫^�E=ź�	K����7��6�I���Iѱ����ѓU�N�nfIb:s-"*ZN�|�,`�sP����dYS�����Tށ�2����B��^NٟT6�G���q�p�W$��ɓ2{~v;&����(`<�+������/��S;���2$`��մ9
����w]H���g��$~��*îtI8IC�>�A|T|wR�=|/ru�ؗ�-��o�U�G��d��wXC%*�f�2"�P�}r�]nٴ�M��e\��{{IŖ�f��=;�c��g&8|6c.x�u ��["�yJ����8��?3�:۸Hxm"�ɤM{���J@��s������Rw��*��AAo��íߠ�b�N��^pJcF�?���Xp�K��U�֏3��c8B	�o��>�35;�o3��8��q?X��J��Q�).Ԝ��t�KEvD4��Zr�&h0�ǈm0��aZ��'^� �Z~_MKB;�?�+���S�: �
ה��9E�ky�9���;�:��U��ld�6��өJ��K��UZ����U��	�{ùt?��-�,��3Ú��}�Ita��S�B�QP.W��=�L�=V��Y*�����V�,,�7r�  �xHE�W��B��7��Ae�F���-��<����+�UH�/�hl�|
��\rg�;5���mh���J�e9d,�M{P��ua߷D��Xa!UB�{n���k�jK�Ѧbbb9.Ʒ�ɒ�;U�/8�G�s>�}H �9pH��i{�a���*؇,�x�ҽ9��
�-�2�n��&���.&�W)�e��]ej������+�L��M�!?\�G\#�gAO$B�>JM�OE3Mn�r[�:�n���\�3�X��!����Ȗ1r��p��)m��ua���~ʄ�� �bs1�f*|�pt⃚�.~v�&-�&��o"�,`QH�?����@�_��ʭ)����!��{Ǩ�sn���<�qԿ;{��栚�=�~u�pfa�і嗸�v�}t�w3da%Ӆ�Қ�%�sWqI������Ǭy��[]� !B5�Ϛu���Y����=g _����
�����#.lj��opTt���L9\���[-ziO�mۖ�N��J&~0����Ćg�q�@��S�J��d�1�,�u�i�c��*����6���/�z�=�e���n�A�~'1�!9�ߐA쎧�<t@0b�IJ����G���",=�%2�~��� �:�,�����ZX�1� Ym�<I�����=?�-��u���5� dD�4���`^_�3��Q[.HHc#��c0o���=r8�/���69'
���2lT�׿��	(m��E f�Dp�_ƈc �>� Z�� FU�'ǿ�+^��O��B�	.z�gU��/�����q��6
�o
m�c�H�|�u�����.��mz��9�Ķ��`n�G��� �'�a������0�c4��Z�%f+���F�W���27�z�5!d���U#I�~�l\���Cx�?Nu� D�f��}��UM���{�ɾlU,�n'��n�!z�PF�Sv�e����ĵ�\ȕW��
��o�.%g�V,w~qe�Gb#7���*�Ms�mNQ���,�H��k������o��$ ".&k �[�dMupf�	W�A��Ŝ�P=~��6�93R=>�)�?�a.P�u��=���`����`�̎a��Ű��3�7�d���Dݞ�K4�hq�d�)������?"�9+qs����D���ݛ��Z�5b�������@{`��NZ�}T^�"���`xE��QuqM������]e�v��h/羽�r8�fZ;"�b[l�#i�~l���')<NM�Iy&�U�����|ɠ��+/Q$��:��GI\�K��_��t��:��%V�	tۧ(����`����=���jI�m�
.%7ZQ$
!�W�oژc{��H$�\�e�o��Y��$'I�A���� #�H��=��y�$*�Z�7���n �����n���(�y�}�ݞ����L]���M� ��g�(���u<Ļ�n���~��E���)9��L|��Y��z4� O=b����1�9�2���S�Om:�s�����2�D>r�'�_ԫ� [���I��~J(2lyx��	ۓ�ܵ� x5S��AFP�8j�[�����\q��`2S�Bӽ	8�n��Jt�|z�_�UyD=����ěOJ�eC�N����1�������?4�5��"w��d�G)�7�}wA�K�pA;����D&y\���{�g ������it�\ʑ�������*gx_���,T҂�Ͽ�vϑMfV���ܑf�9��t�LT��V�C�5�j����s���)-#�nуs랝�O���'��-�WĒ����K�}q����.�ך_�d#�{��%2al���#��s��9����@���;بH/�q'�y;�nv*r{�K�8�1�h�K	^����͘�N�aQ�O�*( -ݧ.Q�c("D{��ş���Pp��:Ҕ�*��"���;	�&�u�e?���P�ˁǑ���"�����v�x ̓�f8���Y�y�vk��͚
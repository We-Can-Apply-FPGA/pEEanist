��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n�W�5��l9�p�9�r2N��t��%�Xm6�L_.^��ed�teQ �*hVp���%���+��U�@_�>���O?Ic�W��%2��U@��eW�wb��Q �J�r;Y�"�4���
e9����*��5��uM�é��t+PtI`�u��w�K�l�s﮹�i�x�{����|Q���=y����m����`����O%&q��џ^Y�V��������0��}X�b�b#T9��?g:��� ��{�:5Q���I����ѫ�Zm����	RϦ�B�E�;�R�
���0��.?��u�&�6��鵀�,�k�@fw,�wn��k0:��@���wӠ/��9}����@��jEݷ	W�C#�ښ��M^����j��*P=ވ~�`;�0�<0KMph��0�'=��M�a�B��ZȦ|t_Qx���3��]�>ek�$u�����T�ǯ�a4)$��zI�g���z����$��+��0>V�V�SgM�)�Ϡ/������ ,��Dwoج՝y|m�v��{!����k	���iJ��;x)�N�N$�|��*.�[�̈́�\Ƃ��a��BFl$��3'��P#Sܗ7#g��)�\�%Aб:�Suhx���;a����JZ�.������<'�o�ʢ
� �1I]_,׈��+2h#��"hUӗ/g��~���zk��E���˶y�!]�3�������}��,=�$[N�Ë\��d�?i��a3�d�ӨAgQ�F����T�	.*:�d��!��)S������ù��-�����z�6��&����P�t�d��p�G�Ig��֚}����ۯ~�m|�x�ud�/��U��y;�����a����9e����U��� �>r�'�^4��v:���Ʋ	���[ҡnR9��CCs�cHɷM(��{Hc�Aa�mMfhѲ�8��~�z����I��>;_>zj���s���X��ݾ�h�&|V�]����)^��,.�aY���Zp9����*^>��,؎��[-�9m&��ݒ9��n&�����_�oX揥��Cw&+���Bs����u�j���_�q�c��,�6����~xӑ���o��VC�1E'�vlh�}HN�u����s���p-]p�{��s��Y����7'T��F��WWx׀Ku�7�R������|�NO���I5��ؽ���o��p���$�<W,��v<Ȅ�#I���y	i`���_���p���ڭ���+r�3e��:����<�pM��Q�䕒�3�u��I��:KX8���0\*υ�d���L��Ku�MY	����ő�ʗ�ς���*Z9#�1Y����@;+��NB56\PC�h��MY�����QAO��I��{|�����V�U���L�?ݯ�eqK���9fi~j�/g^*%sTC	Ӻ_o�*j�Ӓ��C>��Pi�/�UN.Y>x3orz�G�ү�|+�g��1��8I�A��?�2�}�~������"�!o=���K�co���0���ܥ\��I�|#�͍!ۅ/�b_�b'�a@��V�P� [�x�?h�������pj K��-5�H�js ���_ȣ�aU�̯^9;���z��PW�c�N��6D�D�dНC�K��;��b�Y�:#x!N��en36���������	+�\lnG���/3)�ӡ�(Ň(���hF��M���C�/�[�mh��^������P�_!0�����xo�R�N���xZ��XC�3�����E�gPԘ�O��I�{�� /T<�8��2+�f}�염�L�Ec���0��=�?>musT<����]��-���ъ�����QR)����M)r{����2a�F=���#�"��ט�^��o&���l�)_���Y�6|M�;�;����ܜ����jbtY{Tt*��6@gP�;v1��v�#��g#��V�ӀD�,97(۴G}��Fv	~��F�N����jzGU%��N~*�G籛�+����id�̛���X�$�[ʀ�t���/ڀ50?� ��;γ�&�X}���z����Y'�����_��"ë=2%�b9�݀��|"J�\PH���<t�/���5B�bi�Ne����ɬC�2�2�衤i��j�".�g~K���-���h�0�� ��ܲ�z3d2c�wQN�l��j�4N�i ��W9��P^l�����k�%�#��~�- ����cͺ�s��w�����e(���]�#̛�E��giA��OH[�=g�����X-�k�ҽ�$���8����$�Fx�K��,1��6�v	{t9��%���c��!f�Z��0�����#:S�i��\l*��)!��ǳ��w�7@�^�ִ��4�ؼ�C���ڡIi׃��Z���q ^8�F&s�UR]Ҧ����#؂Ʀ�6��ߠ\R���h��W���m�8s��a����\�r����S8fDiC�zqL���(��Zƭ�|7��4��c�SJ7�.��XS�ㄟ�����:�p� �7/׬�w쏑_L�)�{��&������^(��|�C�T�n*���L��(Dn�Z�+m�婻'>�R��xbP�%Q�ߦYNڦ�[��"�9�E���#NkC��N䔕�N��֎�+����������E2Ú��f5z�Eu,r�ۣ��أla;gHCh�B|O�S�bWp���&�Y��P@"E��� g��@�-����A$�� �|�sx���E��Es,�r�$�*$6D�]�ȝ�t������c܏��x5��~mv��F ���9-�9��5�e5��\vf?�D���1��e-���8E�WѠeM2�"�k#�k,����3����x~�jH�6-����Kp�_x�Xw��|; ��}�3]��/�od�g�34�+U��Mu�J��p�nAǁ�ߣH��{#��)Һh7j3�W~>ςMݾgz�^�r�q�	.�_��mi>��d����u���ɰ�]Ӿ��h�q�<��_5_RQ� |�I��6w�����x�z ӣ\2J'H�e٥ !��,1B�1���@�/�fY��n�)2ҡ] 1
�j&Haռ��ȯL���WM��<8�r| �
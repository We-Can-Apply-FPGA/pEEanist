��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��`Ղ���0<a6B��(I�izr��6����,��_��M�:��&�PH���da[��a���V��z��#��bV�#~Z�T�����K���]��v�Ÿ����e�Ǐ�U�F����XPd�}�4T���|�������~"�l�A�]^^R�2.���1ח��:bZ����Q�E/4:�He��"`�XM���xǑ�/��(^H��v6�j��2��F�爴���9�2��y��\�Ob�w��Ne`ӷSK�z�41B���٩d#�*����]�o�܇u1@bMJ�L��2��]u�:#�!̘��*|Q���24����k�)a+��upg�9"�bl@Α�z�y,���q4ꊙ�N��Ͼ{U/�v`& �1�|��P�4�YOZ�t���U�#�]YW���ͱ�0(��r�j"E5�+���3��C'Mf���Fn�:ƨ�����%YnC�g�{m�l��|&|H�&f�:^?m�ʗ�-�ϋ��L��:<��l��W���D�G��m��HB��鋦�uH�bt����hD{���	��yS���ʺ{�|}��`GBB�q�QY�!hg;D9��l���O��W�ܷB����Fsbj\;}�����>	ɤ�b�8��T�/��{;`;�,�� H`�ݡr�m� ��%�_@	b-x�v�����Y���uJr��hM�U
<�#  ��T!����\",��PwX `��J@�o�ľ �H���=����K�U@�;1V0�ٺ�Ҷ`�/�6�͎{O�p+�U���Ϗ�=���J:X�g/� A�+5�@�L��D<*<&0����yTOk�M��#98��Q4���I9�g���!(����ޓj�mR�Nr�R!�W�}�1�7��|դ�(�ݩ���$kJ:�M���%"BDfW0�
L�`J�ps�����՟��e�qs��ƚev�~q ��5�P��%Kq�c%��|�����:}�En�.ޖ�[*|N�K�3�Yg0���譈Ӕ͆�a���O=Tq�W���Sp!
����-cO���R]=0 ��e���fiZ�v<��sG��jT��Ԣ2�@n��\��Ec���%�$3�l��8.?�S��l>2e���`~�p�!���5��pQ�K= N�* �1ɠ�'���7�M��7=����\R�s���~�e4�	�w���iZ{�n<�3�%j.�E�E��\�4��x0��<f���=��G�߄��5h�n�4�<��gp�Fl�ކ1���K���;K��ɦ��v޿F�"Яi�e�R!%�yv npal�>;���P�I�z��Bn�4h�w �M!��D�]>��2԰����k����	����!�����Ͽ��~������w�}Y��8��a�����k����<C$@c �ך�[�nS�y �޷N<imƲ!�*�<�M�.�.N���^V��d$v=�AfH��:S����b`��������}}"�{��)��x��

W&����Kw�U<@_]���h���	9j1w��z:�c8�L�(���ۗ�|8�¨?�Kx�2��a����ӕ8 0tG�j/�ĥ�����l{���H)-���z��[hZ�[Ao����{���6��A��P/�`"�}�x�u��'J�k��j���&mwI/��n~e���ވ��P��u}�\��F����"?�*��qG��j0#�Each�����&�Z���YJE{deT��c�6in���_
W[n��]��1=9'�R����!t`/&����YT�bN��G�j ��_#}�����}�7�O����r�P�nGk�̼�,!t>���a�}-Qp�ϙ�JOy�rU�S��r���w���:��5������k���w� ΁��I�Ûь���jG	�����1!f9|����.��'���F����+�9_���@�׳��ٰk��_d%�ɽ�R�9@�"�]�ְ��G�#2�_�@�.�T)�rCZ�;˘3�&B���~^|�����k���i2�ٹ�F��y�i�N˫���T���՜����.k�9�N<��v-��	��/��Ų2ȔF���l@���E�d]H��]W�v���4 ր!l2z#��?B�TN�a�q'�,�y��1�*��S��0�B�b���@�6�+-Ac�ɦ� *8��<OҮ �����U�(���>q~���g������h����Fr�#Ey�΂�Z��L*�}�_I��/;���Ҍ[�
�g���I���(ݥ����>��,�7��5=̥�ء��Ҧ�����Me3k٥0hW.Kl3}SQ�~mu�<�K��a���q�õ+m�Q��:{�[��D�V r=<���U�D�0���� ���[����ɂW�.-FA�}�E�'�0����g�I��R�����c6���� �S��;��0�X�=�;��Sz�z_�=$}�耎|Z�T������������1��=�ȍw46 �O�6@g��ŢQ%��������3�S��e������E�\5���@(Vl�aZA��NH��/)|����4����q��ӛ �̿��єG%篊��)�2������l�_N+���F�N�Cp<>��ħQ#���ΐ���3�����BC)r��R�zi:Í� �>-�t`�<$�>�9��iW�,[0؄
���
�q���0�,JV�}tL�-�DC8�-9�q6%�����'�U��&�M��2���"W5����n�����:fX��hyh� )�S�O�+�9�?p��̜�~e�
_�E'��dz��7��P{I��֨�Q�@ۥ;�1����lt�� ��HV��p�0x����lJ��*v��� �3�Tu0�"ۥ�`=�k�ij����H��.<i��B���T��F���'�k��1���l��)yEI�0�[�&��"7F*������˵N���b�R|��_p�=�6��r�J���Qm��[Q>�)g���`=8?��S������������愫�s���W�.ʱ��Gq휸���U�AEP&����xcԏ�ɘLa�iB<�C�x�}�J!�KQ�|/�c�*��Q��� ,���N����7V������BŹ�ݹ�>2�٘�F׋���8[��*�1&L1O;�3*�+��+.X'g?خU���frq�1����Tg��ux=��ƃ���<�K(�.�UhP�'O���+�Z�S5�7v|ٝ2c����zMȪ�q�'a��:����M;�^�UtL��<T�K2�e˻5�Ua.Ңg,����Q�*6\��5�K`uJ��P�e1��J��*u��{�}�3G�hֳ�L�-�J�R#>��֏��[��ȴ[�����lQY"P�|T6
>����:�~��t��%�6�f�\feݛ�,�5�&47i�{�������?I���~��������|J�'5i4�En��h�eȩ�ټ���i=�(T�����y`�]}�θ,j8��X�F�|	��ɌxQο�>���;N:0s'j�h?n�ֱV*/�0V�q�'bu������C��U�����r9�	e�L�K[�J�4��˄��gbT���Vg��XĀMu$�|պ��D G�c�ne�C������Ng�r����?��(Ȉ�0����c�R�^C�A(��#����Hi�(���J`Y�v���et+�	>2�. X���aWoZfI���	�ʌ�7T+ �y0�f��VAIH!���&']�Y�n��}G9F_#�>�ã��%p­ �J[�)#���do����ox留�1�J�ˑ��3q�ק� ܸ�S�6���e�t^��R!{P�`��ʺ��ki=���*�E��#�������#���� �n?5y��9�+���7�hs\?6ćߡ+s��ܑ��������"��c��Z���E��H�ne�ۮ��L#�Ň�S1I��ߩz���:Cq����6iF��TL������!�	���r�)S���u������)㾰�w����78R);�?�kϝ b��ڒ����e��5���GN��M�N{�?w�{�����h&����� zW0e��D���7�q�&7V;R���;G��v�ƭN�l�&�x�KT�q�!�P���x=q0���]�\hz�^�Ԍ�����U�����.T6�A����s�����G�j� %g �)��n�r���a��D�@U��
qb�c��ĥ@��8�LOmp!h6�̻q�
�����at�?��P��ZiJ�	;�D�1����yx"j@�;G�����`(��
2N�e��+M��A"l8TFWd^[���a�u�2��Pg'kJg��u�9�`Ci��ق�Vت�ZM�.;a,c���ō�qm"�m���E�[s�+�:gWl�TS�]O�y��*�`��F��	Us���\��������(��N�W��O���8a�ӝ�u�����G��e��2�wݧ:�<T�Gy,�r�C7�k���Rq{/�i2N�@YF��t$�G�Pĕ�"�A��vch�z5mL��U�&�T�GG���e40�Yk&~��I�����1�?K;�#�9k(��z��T����N��!�iԶk�����Gc�E��8�|�
�sYY����̛=C�U�H�!����$5ƨϸ����������tX�QᾩF��:XJ��ݚ-��$&Y_�u�ָg���� �Hz엾<��`�8½�'v-:EW�-=	'2eσX�����Ū&.�d�U_S�.��Ĉ����Fg�'�P�w*�MAn�1��Ӡ�yE>4	���\yO�aA�lQ��c+��G4��ؼ<�чa�rs�Rꢆ=�}C����zt�aO�QS0�`P-�0����JhK�cЃ���h�;��цF3�ue�O,�gB�Z�&�N�ɬ�YhJR&O,,\J�����欌{��8ll���]:)�`�ft1'��8ܷ'�?lN�Be�Z���[�	�����'�@P�hs�¾�H/h���w��j�9�=7�m��_���$�x����9
���\�A!�L��{���a�9>
)��E$�
�c5��r�Ӻz�(�+צ���i��֪/���6=g�~o'ק����+<�$1��%���tʥ�V'�r�`��M9H�>�1��%)r���je�-_�����p���j��w���@��LjL��Q*#ϗ���h�q���b�<�s���8�U�m���\�BX#N��/U�* .�bV����jX����"e�
43�,���<�pH�E]{ ���6�x�Os���w}��l7L��&�D���"Wz��Zc+9?GB�byj�}�;�������̜5^�M�y�/5<jp����ۥ����s&�^�3n�Jۧu�ĩ����X� MZ�F^�]��� ��H?�H]L�G�Qq ��d
oW��[�Lxޤ�=�y�
�����tƨ�����B����A%֬�jv��4�0�S�o,�٢Dɔ1:/s*�(�+���I��9NZX��6�76�iW}��xu����u�~�^9��b	�g������3�k�r�q2�p�O�T%�"���LԘـ8��L�f��z�q8����<}��w�'�)~{ I�*��u�KG'����
�|��6���Q���ܤ �B�7��컟o�*��K�~�Ȇ�ُ>e���>�Ԁ���c��!6�rw����M3�)��]�[c��Ǽȓ	v�x"��a�C���V��#.2k��;�!w�,j5��>}�+Q9yr�y��$�ER�!�#�ᚚl��Q��oݦ�e�>��k�	ͮ,؝�u�ۊ[�����V���.J�V�����_D�~�[�@����@�0=�L �5���P�E������>lkG>�$�^?���10�g#N����kv�k�?�������fx��O��(	t4쾻l�X�C�x$t�`i斺F��ic=u��[�Ă���!�T��n@��6��n��ЎIԇ�t ��M�>M�f����g�+�ih���f������:��������?�y��ra���бv�Gn%=�v?�������=���yJ��x;�FK�$�.en�z!�Hҏ5dx����K��
O�U�mض�|+L1�E4IW�Tfo{�.�഼ڧ�,��R�[M��"�N��˟@�OGB�N�	�%�?f�*ƒ��uVٰEG�?9f�l�4b��)H�O�C>�Cv�k�.?�0o��F�~/�A���knyjO�K�k�ԯX��w֬��p*�jƲ����YPƘ��[����B����}�O�x�:iT���L�ee{�����DNN��~}��a9��ٮ��S��e���:4��-�`��x#&9��B�����4}�¹?4p�����E�L}��{*�d��*�֤�+Iuʆ�>�����T\LNi�Q5*�j�J
%-�ÎVoVwHN��'�3nx����+����\�,n�w�_+hn���z�X4��}�Fù�!�<����������NMH�۹���@��r�_�b��z�Z�8��CZ�n,S}RQ��sNs�?��*�������'qu�I�������5$ �.��9~�yb����U���A/�Z>����C@�m*L�SU��;����t ��/4&`���������Wd�N�7��1�r���Ĵ�/+������J����{�1�j3Sn˹D��V�E5ir��1]��������܈��� ���:�m�:=�>��J�X��z��_T\��O�8V��q��4� ��Id��,BnT����4k�A�])!AUّ,,�-,����kÐ��k�R��&�&�А�Is�A�Ǿ�������+ع��BL���>h.��W�a���t7��n�'�PN�c�6"�L�����d��[�P��!y�/�3�ڍ�����MA�w^�[���n�Py�at�/�|ǯ�1&�l&cQ+��祡↞��o��aG#�UT���a����6�ٮH�M~�r8�Kx]&���hrI����g��S�ak��������R����[�9��2��
?�"!��Z�1ۥ�l�ɯ�����?E>�8���H;��k�@z�X�]�eZ2����'�4&c�T�H�:?���|A����*
b��p�ф���|�9xmh�BH����UEM&�	��ֆ4'Ղvö�@���^Mn�lv�3lU�<��,���5���<G�dv-9������L��&�k�B�/-af��p*�L"��T]��F-���l�_��f m�mm���e"w�x¿F�� ?�JY��.���^G��.�)8q%P~q�Wg�U��^����q�׫�́m�l<<f�Z�(�)�爽А�ß}3�[E��{� �7^�bN�::���K��s�;�N��C���³h�����.r��D:Z1�.��h�*�A�!�X�zM�Ӎa��[��j+�ՔVpi�q�78� !�§��o1�jK��Vw�A4��Vژ�)�`��23zea�is���F�r��iv��d�7.F;��>���,����4
�M��0�Rs���Z�Wg��x�eIufA�hˣ\^N���V�r"c�y�����\�=u)����9�����7's�wG�0���	�%GyA@d�k��>�L�P�	�Q$��&�����Gr�u�C �$��kƐK.Ɠg�US����l�t��TW�^Pph�Ʀ^yT"$����rT���~�{��IF]g�*�7t�^����û�ʅW/-.K�is�|�u�'\��2 �(�B�u�^Rf\����aFz1�:�����u\��S�|���ʓ,����4,*��g����7�95?A�[����_�񞉝+GuT���b���_�l�AE7��?�?oVV�y��}?�'�oLX���3�:�I��(C���t	#�cX�R���w���L�6mpb+!`�^��)y�{SE�P0|�N1�W�T��};��lw��J�ۗ|�!����^�pZ�틀�]�Μ|+&��&��p*�'��,���4�!�&�"h�]��\� {�H�݅	�:�T��͑a�16Ѵ۔�5���j�U�w�\��,�4�t�MhA[�V��V��b�RT��Gɿ������#���Wn�ڣR`TJ�2�:��۫`�{�-��}Ӌ� �����*?A��5�L�g�p �6���ٴ�|�
�fJ���,b!x���W�<�ջ
�uQ�����W�n�>B�?��]�an�M#����/5N��hWN���"q�xo7J��
j�W�f
77�>ztf�}$8M�ipe��õ���C�����<��a�ڨ��f\+��!�GM�у@)�:����~�G���Aai� Nth^7���G�@�n�|9�M�'���NUA6a����˷��1Go��[4������`ֹ�J,��ˎ���J��:E�[���E�w����b����+�
�n�����<~�H�f���<R�C:v������	��������nm�Uy�&ъ�պ/U*@[͝=�/���;�P�9U@hs�<F���~$�:��[e������PZ<��y�h���<J�+��\���kC7�0|��Yz��,���Qjk���G��z�9_��Б�z3��)u��m���*�o!qXW+��a/�Y� �o���
�Ɯ⫾�~TIn�#RL��d����2��[e��%̷=$S�Fp\�d�Z��8e�S��0FF�f�龀��^��̾4̓pI�n{WGbZXv��pĢ�`�W�{�Fҧ��Ȋ�V���x	����<�4Km��o�3���EfmҷQ�����d<��Ћ��s�.���(0C0����\{�\X�WX���4`�+�G����60����o p�<eU;�2�
8����6?��$������oBT��),Bm�/c�;��66�N�9xҡ\~HJM5�ʹ���������m���į �F��K��_��5�F(`� ws� \4�Jݥ��*�B��J�nh�B��b��9G� :��8���ֱf�v� �=����8v8!��ޢ���g՝���^��R�/�g�E���8�������3������`�[���P�ɿ��Q���Y:���tyrC��׏�$��|2'����Z�Lٸ+�v:�4X���*D�,�k������;)��%��-��e��1�O����Ԋ�wWZ4&ɜ{S�xZ:5}q��您ƾ���b�|�kQ` l�ҋ��-9Z.~JJ�_i�j��!3�W�A������&���t&*!���[�=V5qʭ�@���?���"�DPs��WS���@Xg���w7Hn��d㶄p��c���H6X*��"�z����׫
�l�ӏ֭2�^�"�%ܚ�B�=i�8�����sD���XR�cמK�tSȚ�䣈J��d�L~N;,�|��[W*q����cb����D���b��	����#lm,޴���k�4J���T�{c�#Q����٫ɐ�+#��Uh�e�t�{�z��\V.f� 6B��_�X�� �Y�7OE��q�s| ��'��l��������eu}���\���з�7HGm7Wo޼`*��.����=���*�ߤu�V�w��Df܄�׆D�q
��0�	g�&td?�1�tA2��՝@�BЈ��N9�P��cm��Ǎqr�~X��_���3%��0���� pr*ٚ�Xd�Ah������O_^`Y�=��;j�lt������� �t��,ŵ�%��:O�܏�C�:��������r�OU�.4F�ȶ*����y�S�}��9!?��L�)4,N�87�<�U豛�K�0�Je��\��r	�����$�P��v�X���z�^��;���_�w9�%��Q�=�ٌO"¯�̠9�g�*�W�b]��mqŋ�R�hi��'��v�]UIT�t�I7V2�)^�K^�G�{�A��a���U�@�ݚx���aև]�i6��<_F��ŀ$a�9t�><��9���>o3jbħw��3�@�Es��a�P� �j'P|� ���˹��qiB0�<�*X�OS���T{4��-�,ս6#���)AlL�@j�j��x�Q�h�$vsă#}h�������d�փ��l�YV��\��_kO���=���q@���\��}�����ѻ�	jX���:w�%�H��nQ|m[����0i�C�@'�47�F*��dB�5���u<����Ϡ��Mh��\�3�!��z7��&�y/SB`���|�
ds��ZњQ�mj��\��<�dif��
%��"��I���`ZB��UP�O��8[�����O{�1^H�/�֧�;L��-��re�M|�u�gc��RrpaY�,S��ϕ��p} K�ݞyX��_@�ŧ_�[M����Bd��d��d���Y����s<rb�ē����u&g&�ԇ��]�&�uj��s<f�})�*L�rfG��,���[-+o�.�iR�}'�x!�T� َZ!m���*�|�oȿ��
=���<�	x��:�)5>'��{��T��Y�=���?�1-��e��f*�O�ñ��ca���2��AL�6���*�PӸ�y<��u'
��g�pn�'Mj;L	�/�;�#�Ԛe �@�%����}_�jUo����p���Ƒ�
�ά	��ٱ��:*�`�{�׈~����.����E�%��ѫ&g�>1 /&��
n:�RMs��&.����*���m�Ffl�;+�Z�S��@q�������T��+�����Vx��Xuۯ�Er~�b��̇_��>��d���s����f6(������@.3�/R_5N7��V-*Q�+Е��efa���D[��+�Q�7�a,���vi2�;�U&�����đ]<a�ymş�5��r�S�Be�G�3ڌ�] �$��A�8�S�>D*ncl����z����&)<��k�����ɣ�+(���m,�|z����/���Τk���p[�v�A�Gʉ_j�9J�4~�`:�L)��)D	Z���J	p>�V���3�Cr�{mɈ�Dw�J5P��,�
�<��#��TӼ�~�� �]I�Tq���&��'[�m�DkK��2*�}]-�N��4��&�w�3��e@d�ܤ�߱�J 4?�����Y\�r�U�\�c����@���5O����I|������bW$�7l�m位d�=7n���6*f���\��ԗ�a: Q��_y���-�`!��a�)�U.v�;�ZO�|�qf�p[W�#:1�hC[Yets"9͏�b@�(�ڦ7�'M?\`��E����"Z38�����l�����(�FܒIN�5�Dz�;��a�d@M�ӋL��g��t�	x��8�D��yQ����3wjG���|�;�ڮ��L:�! ��4���S�!�u|h��?�3�G��,xe���`�9Q�n�bX�s�+dc��%q����V�}<�81 q�&�M��~i��o���qT���>�X��Y���7���Sy��4�Pӈ�����*�pȺg��r=Z���ĕO������`8�,�����O�O���ʊRqؖ��`����і5=��\fo�<a�>&��>:'b\xX�Q��J�ɾ��)��	�ђZ{;�!n��ۭ���=��˒b�R�Х����{�9��*�����b�Zl���_9�P}K=�=�O�l��]h�bV�*����D-��!67�e��`s͟� ���q ��� ���̐����Վ�XK���UQu����MF�ӛ�"Әf���g��f!Ve*T�u}��od�^�=�wLJ"�	o���,�e�ua�A��k�P�u���Z�f���p����w�H������@S��̅�{�)�E1�Ņ��Ӯ��El>�jޣ��L�ׂ��
L��z��M���E%�� �Y;�Pr��i������va�����JJʹl�g��I�3�g;!���'}��:GD��r���d׫@ޜB�k*ad�|ۉA>1'�����X��8 �WE���QC��Q$�;zJ6�76�;HK �v'�|���d�W\�}P�]$��Di�=���-Ї�;ov�XB�'�~̷�:iU��BZ��
�#}qw�L}~��9�4�K��?�"�x@;���.;�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n�z���Ͽˡh��ȳ������E"J��ʼ�U��;Z �ԙGa퐁�o�S�`giDh74|%�q�/|�N���E�N7y��x=w�s�6#*�k��9ɞt���'Y�dQ��6�)ʶ�IL`~����I��x2'tr��O�h5G�Q������!|���ak�
�}�
�i�c��.�)��Gr��G/A���.Ӆ[
+��B :����c�F��`l�f�+���}°�A��"sޓ`���|�5�46&��L �~��ds�`�s�מ5��_����v`m��!`vw"���f����m��tz��K�����AE�<�E��|���f��*��G ���:�J��b{�I*�9k(ݩe�;���s!B�uN�i��a�#eV��E��g���`F�����kI�����<�/����+P�b�Qd.��^�s֜g�x��"b�S�"�T5�E�X_���5k�г )ί��,�?��f6aЂ�d���Ry@O+�7�<7D0�6H�މ��Gm"����D
L>��1ޤ�a��ѵ��3�ln�a�W��hEb�{�j�1���G/Xp���.0bh�Q�����b��?�{�TDӑ���;+o���J������E)����F}�WI]W�M�8��㰟�C�.x���~��T$��k�� �Kzj������WA�
d��C%jJӠ	X`s�����,� �nU�`G�>Cx3LF����(�a|�$��h��s����d~:\w�O�sX�ڢ�����3h�rÚ_�a�97�dAc(;wm����,��B��C�'W`k��ǃcJ�/&Z.��g����N�J=Z�~t�s� ��=%DO�
��x�@M����I,��c���t�t ��n��>��i��#J"��z�a���}؝��	g��Di�}.��:�弛`/���;>���)n�6@㟾��9�³����O8_�(oo�nV�.eB�H̨K�F�<B=��6�tux���d�]GW�M�F�U>�%7�h����+���L�xvS
��'nP�b���%AD$�V����!Esξ�2?��5���������F��TȪD���r5/"~�cq�&4��j
����.s�c�*�G�AD����,pn'P4��@���=�?�d�B@�YFF��oA��D@5u��(�����l�a�n`�������Ϣ��4u�J��Xk� ��h-�HYv@�]�mp�7����(V7����-o����礘�b��0X�d:"��P߉U.�	at����%���a[�-�U���.J�P�q����7zˡ�h����Q=�y���(o�\Gg�!h�Ԉ-�%,ݳ�9s��оT��r^ͺs\���E*��[�v��}x�e���6���o��eM"
y2� ]R�l�#wH��-�q��:U��v���?	M����Dt!M��2Ό)9�m2��C}#�-9�2P}���G�p$��l��X�
5�n�e����f( a'T��P�Av�''� \��4�U��X��$IMnS'�������S���й� W��`j#(>4?��ԁXe�yqA��Ҳ>���\�aR�(̐�Q�"������^$M�	�q]:��=�5���Ĉ}���hEg�:5�Y����&ϙS���u!���$��gHp�Ig÷��P��:5Y��VRu~��9�E�ԕ&�����+�p|����cY�y���:}�?��!��㕅X�M��n��!��۰ѣ�+c�L���-[�bA'Z�qn�ŷu9�h��h��+�X<ǅ�t(�u :�9����f�W⴦szR[��|9ٚ}�f���� �]W��1��J�F��,PK6�3���t��9��8:��~�á�z��x��8J��5%I9�8��wө9_o�FY�Y��+���kCW6A�\)X�Hϣ�X�\Sq+_!�TM�"�B׌����~W�
�'��Ͼ��s:�~Y���\���\|ͻt��[op���N<�(��u��p5��G�n��a
���ĽՋ��K��a�1��������(�m+ՏY�{��Ɨޭ �8998�Y�N���z�s~M4L��+�e/vS�ZP�,�#��"R�Ŭ�1$�{67F�zo�j�� �6��~�$��2?�,��r\�_�'����p�¾b���AU��6'����NN�����H�%��ߊq3d#"��M���[SE��ahڨ�x<;ʄ�>�H8I�}k��&x��^Zu�3~h� _�����R�q˧��t�ŵ�6t���;L���u�	E��Xm<{�d�$� t�M�Ǯ-��M���RR'+:S2���\!+-7�����o�o�l��Q�M�Q�Q���sa��Un��x�)O�z��3j�������v��{�C�4*``�AL.ݙ;�������b	G��+7|1tC��Dly�2*z���{7n���@@xsJ,���?j�bQ7������.D֧����9�qY��dS�dâ~ t����Ca]�7u��$~�Hq��`j��ӰB��2�H���c��}�&'�����?�OK܅E���̤VQM�l��G�03v��� ��
[�j6h	��=���SM�/����H����<�#K^��\�~�ƕ{�d;w��L�G��u���z�T1�ҳ�q�R_==�_�R4���f��l��) a`~F8��/k�Ax)��K�i��K]!3�'��{��������{�����q/n�3�@K�Fo	�Au�Z���I^dY��B�1��i�\?��Ub_)T�K1�1l3�xR-�}p�<�痘2�s���=J�x�� ��k�|ٍynO��>�Q8��hs���8,1^ix��@Mߥ��l��$+����B��%P�k�2m��ݜ���M�Zx�.�\�PI)?,:�(`�"E�EaZ_.�)���7e������o����f�V\�5A�u3}�j���p��߀�Z�6��R;������EO��;&�����k�]�eOI]�ī��N�[�JT>��J.W�1s*��?k�1w�����4��i��*\t��źNS7]��v]DGm��%n�9"2ϱ`�����>r�*���`��I�R;�t�e9�ۤ^���l	��v��>rTEp�s`;�u���Iwk�`�+�_n\��Q���d0�	cS��z�w�x��� ^6QH�-/��J���RB��qh%c_��֥��.�"�5��l�dm���_�L֐����K��T�>�e���#�kڶ6%��ݼ�5��q�!z�g2�p{+��0\���ڮ"}� ���?�F?�y�>=�x[�øe ����ιY�-�5�N���9�'�M,����8��~gp��>��\(N�dٷyH=Ṉ=l=D�,������|VW#i 5ޛ)d��{��N�q_Η�;�Xr_3�e�_�n����܂W�YuKz�0�l�%��DY�/{Cusz��c;~��=Q+��G�[N� �,����u=�� �l�_'�r�~����&�:i�UB�������}�A�cy���)�nx�QT\��\ˎo^w�6��*)��:FIS�����/�`9Iu� ��<f�D��Z��5NG�e��ve��'���9�ì��X�)�X2	�����,f�ڱ�i	Yi֫R��mu�Jd6q��r<�$/ǆX$�<��Ž����Cb�C�ܱ���o��4Z~1�][�c��f�+L*:�s֯�a��h����*�e�%�2�A�}�8��/-q(��Ǉ���;�(6,��E���[�JB~��-�=G�DO����L�_�xv���̀�툀���F$P�"7�(�z����R͉$F�϶',��,���U�0n�	T�^�δ>8GK�0�@�v(�e��xl%�Lvݏ���s�w'���hM3w'���g���ߵx�"���I������o�P��$�J)�jf~��Y��I���&�3�kz9�(V�~c�dq뺎u�Z.-	3?h��W�"[ ʦ.�J�{��kp"L�8����G���OY	q�,>��tRK�Ic�贠ѫ�Y�O�p�����@�33-�Tp��{Z>+=!��� ���6@�{�.�Z�I�+6'���� 蝹z�tL�.rO<R0�W�Tw���Ғ�*m��$n�*�2N2�v��ϧ^5�4+Y�k;�g�l�a9>�!�5�W��F��"ݥ؅��e�D�zݾTq�>YL'	=Q5YK��y�\
��.�	�ۭ�_ҏ �a�(��0��w{�h��9��<u����o6�;���ɔ�eO�$� �32pᎆ&c{����ЋعQ2-�PPx�-t�6��8��ܦ�ͽ��V�o�W�+^m]�t���m��=��N�Q�}D������(3��8V���ݡ�:��O%n��Ӏcr�?4�gf�%�|�N��m�e��F��M��)l-�v;r>�� Z�	� �3��B��w9�q�j�&�f�H�v55m���|�!��d�n ��S����Z���1@�7��@G�b"c�3(NMK}8�\�	K�(g����цy/�s��F���
��eq��:�>�S�<S�SP������Ք���۔	0{�tՐ�n��7y�P��$t5,xG�>dA&��K�I �v�O/�\'6�����z]��C��B���6ܖ7��z-�x�m�֓�����2n��Յ�U��kmd<w�R�ᓪq4�m��x:f�yށ̘i�gɎ��OCF���_�	w�;��Ǖp�u)��'�S��V��x����dS(����5H�հ~lxy&9���2S�H�Ju�F�{�}'�@��4ҋV'As}&�ӌW*L�������s�H��#>�=O:CI��M�z���c����)����	 ��Du:U��@���L��n<���M�`:�u�>+A��q����hº�Ml��N�����yB���yϕ�O�� h�->����R�.<T�<5+�������O����^
�I �:�B�JA�%��f�N�kS��L�%O&������ �LPl�@��vJ(�Z)�� ��L�i���G��V,y�D�/�%��PV�f��B�[K俫]y�,
�I5Yt!�X�1�Th_�l-c�[�hP�g7��sO�X��]lv�9�	�������)�S,�����fT����X���bn�:��^�H����n!�N,F189C�����O\�6��a��.�c��4nI�_;d����O����HA��c
���ku���H����~7�9���:�fkC����_������~A���z���A4��
��3I�c���>HӬh�T;�_�|��b�ۊh�����5g��.��¹����	����@5�EK���O�̅A/�]��H�ݐ!R����L��!ϡ�c��H�\�]@T���2�׭:xQ��h�*�WJ�v���W��kc��i�W�ц�ⲙ��X��{gk�#��AV��OC��dH�����,�E8�㾹&c�g"���/��{�Ӓy�7�2ڤ`[gʠ�j�t��-&����s�`�����u�H�Oӄ��ٗ�S'�C5]�^N���	���	�/vn�5f�_���ay\�e���<f�^�ߟ	�8g봉�h����C�Q�=&ozO�K�
&V-�m~�kq_$��[���/r]9l���6���\�v#�F��
>͗��&lXFT4^��-�X-�	q�����S��l
ZN�Ȟ^����]/Ҧ�.KO�h1����8�u�	Ali�<��Ѐ��q�u0���=���;j��XH�6�:¬ݡ��i�� F3R�q<#��*&�`魈ئЯ�5��8�Dl��G�T�Ó����Z�+�/�u�It@VCr^>a��O2��Oa��1*�i�~N�E!ƚ�f. ��d���a��>唭����B�e˵�>eڄ����ze����[������uQ�[q&zse<y?p���Q�0UN�\�hc�otzy�V֧:-��؁:uԝ��ӗ�ڡ5��5x-ۧA��E�e� ��I��������6�U�x�L֜@��-ͱ�cy�^�*�����o��3�w߼���s]-FT>��u0�w�_	g��N���EL��\�	<\'��5�7��"H��cN�hB�w�MnƖ+$��1����j�,��������Y�m�X��RԜ���@8��h[�����h�3N̗����m�|,o�b��nq*�h��;q9)���̽|����_.�"��:�P�$��~l�m'VV�q�G �O�����ێ0"-����hN�z��sԆ�yࣉ��ڮ��Mޗɴ����&�[�n����|�PP�ō|,D�-����M������(l�V��nϵ4K�7���bx�p�r[�ä|�pqK��fV�#E�,��͈=�pNl�5�Rg����I��,�%����|K��Hܐ�/��e�	UQ�1��k������\���ư���.�u8I�h��H��0L�;�7�Kf.	t�2��ܴ��,_;hG�5��=w�&j���2%Ib��4�mL׷Xk�����p�V����<Z���;����2�:h��(L�=͖\3.h��	-t�(�ؙ�������@cv��%2"S%oW)M��q�����#wWŘ��űଉ����v�L�������曧<&�P���I�H�Ò)��W�>�����HtP/xTu�^NFX]GW��������h��d�si�5�,��[�J,�"��FO 2��E ��ꦀZ75&��k��qס�L��1�ć�2M�ۄE�����\�as$Z��+�{����铖o�~���ϱ�:��~���Ln/���x��^��IR�i,4�I xС��a��� M��.+p�2w�q$�L��%��t}J�u��� �[�$��6���K�>&�t�
�1�^�j�f�r����HB���w�±�뵝�L���4��G��N��w�Yd*G�{��&�L%⤊��h��:bL��[��K�a��1��սG5QnX,�Q�5�U�F�/E�72p'�U�����@��o � UZ��%_�t\랭�m�2��)ެ�mV�������p�2 �?���`��������U����G_5v�����
kȉ����:�L�|�J�(��]KS��?f���g�g�ך�9V��.�B��ǳR�FE�
�K�Z�:�J�;�T�Y1!z���39y�\��S����������%)���6�����/��*/�!�%1H�L&�m��.X��?%��i��^a��³jx���؛�˳~8һ�C�8I��I���~��]no��~�ЁM������+�9,r�r�%~r}zF_��d6�H!��c�=?���A�bn����%R��5`-`�� p=/ݾ@A��#���-t%��Ѯ�+� 
&��d�=���EFL�_�υ����P+��Ϋ�tW�w`�=�d��|d�.�q�tiq��EC��L�B�)��>�M�<�!�6+F�O���b��e\�c)5���5����+]�z���M�;�-�a���w��z�b���7�������_75}���u~n���m�3e�ߤb����0�O����>;�]�6wu�Dܒ�� #�mh C�=�O40��_M�в��o�&|3 ��'f�3䗲���U�V~U(���ҸK�>C��w�7��� ͽ^�?J�&�^;\�z=XψK���1#����{%��r��CM�L��^�Z�;�T_9+��e�+R�����?xV<r�ii���O�f3�����i߻�H��ԕsո��/v��Xڶ_�E�bi��`(,�9���Җ��J��|J̀���J���{l��љ&��o�P~6�G�_�m,}�{�xR��*���[����Ӕy�?"�f����+E���u�A�y�F^lh-��4N�`��!TZc��'=�|t5uZ�肄Sh��j�d�"�����ʱ37�T2�r-�{���\�#�v��ծ�8xւ�.[���C��l����#D�ZN~_杪-J�/
�tRߒ}14�G��V賆���t7���X�������@*Z7�J��O�Q6ۂ�6�[�:)Kp�p���npŢqr$BѰ����4?�� jI�R����9��>)E��D�`\���:�V�0�1�Df�?e���˙������[#�Ơ�~��K�JEn����0'�h�:��-q�M��\�x��cH�U��v+g�|�5A)	�'���,���_�v�%"
h�#�(U��o.� L�h��e�����5aX�=��C���-�v��G��%
�!��2g��V��+�ߩ\b�>�$��0�OJ�W:�^���I��2SB��f�:m|$`��L�,�Ӛ=�K@q d�b����00�M�߿����U��I�����{5z��f]G�k'
�����HL��{\�k�0B��*�,����)Tڐ��f�.�x�I��7$�� � V���9
rCH�B�����b��0�������T�!`���4�I�{yc3�a�!�p�4>S�6M���1�z���a:�I5\��)�
�e�_k����oB�� &���c�uF��p����_Z;��,EA�AǪ�к�$��+��穞[�=������:��O��9&B�0t}g��&8�;��n�b6A8�)�+���$�ㄴ��YQaU�9��Z}�a�!�v=��}f�M�aM0�B��-�����Vk+��0;:9�&���۷��mV-W�լz�z֕��%��A^DwX�2c5��l����!)I���r���]fۣ�tGޛW/�wKtao��)~q9*��T��������N�͓�}�p��jbʦ����-�0��<r��%Q���@��x�F��1��[b�)�1�eÑ�.�98j�o���-a��[u��QQq�̀&��p�␙������
*��K�k�w���K�'
���F�4�5��F}���ȫz| ��m$�T�mE��a�����؅*<U�Q/8�����a��ŷu�Q�gl�T�D�+ެ$wY��_}L�a�f|�J��9�䧝����B�;b��ڽ[�r�ᴗ
o������ SZ�����R�SNv +��K��sx[4nQ��IP;���<݌�l��6cw����hQd%LJA���%���G氜rP�У,��-L�QD~��'�v��2�8��o͆�H4>⊞�VGe ���/xF��{���E�1>��$,<������נjU�эEG����Q<�E�����q�Nq��&؅���e�P�ݎH���t�+��)�)j>���a9����{7�?;�*Rt�y�F�hp?�JM0?r[���]����|?Dj�ObR����]�����k�0D�.?�L�)Y@���k�줅�J�:�&n�t��"GTg� �A�#�՘OW�Ynm[��̀~�/��[Ibw���i�`cD= MY��%�h9�/�*c]��"��*Î�<��	%�}�dc�>�Gˍ��L�'o&�ذs@��o;_|���s�2>�����4��Ǥ90��$�8�Fdz�"��
�-0�+�G<��(rr���ʖ����?=*1Oj�FJL���O��,�٪���qJ���8%B,U�q�?����	)�����r�����^]>�$�fv�s#GC5B{.�K���x��V�]���^���~(˝�)~͖�V���2N��vIP����'���xM�pL����<u|��P��X=��Y��%J5k���.�I�\TD d�:�Ⱦ�	��$�^��p�KסiI6�!�;�g:��$K�����f;f�.�ch=��^�Q��%�񟞦�����o��!\��ɯy��dCR�q���������~:��J�O���<'lS�W�A��f����E�b���n�#K5�ʽ����h�LD�l[��R��:��L��먗��d�p0ѣ��j^Fli]FTSQ����w��41X��|q�J���ѝ�ŶO��~�jpr�)�ώ�7������+<<?"sX��;^���qvW
ehW�ҩr�I|�^�35�+yy�:9�ZB1�b�t��Wד)�Ƙ�#���+���@ڒ���r�v�R�A^��|�JMjD��l�ڻ���hࠃh'�	D�.Ǎ�Yi���V�AE{����N���e8@��W�ѶoK��i��{Q�8qȅ�;�
5��&pY�D&����	�n�L��K�F�M�
?f˱
?ZW�����ͥ]�c�y�-
��o�t`�A�1����ΰ)����+g�d؝l��K��͍���E׌����\3u�t��Kv�y����Z&?��G�[�ܠ�2��K�m��M�.�f&�Hkk�Z�����v�d�#:U����}�y�K��Ļ4�CT��-m�;-���Aqh��M+���9Mgp���oϳ>��aላŏ�J?_x�>��7Y]2\��7�En����Z~\?�W�Ui��c��қ��D�1 ���Se�5��H�b�D��n�^@�y�o�!�����+�$("�"1���l��J���XC�����=d�ǐ�qbs�����s�m*��m<�B�T�����ʟ��.��X	g%���&���\ڡ��饚t��d�QQ��O��l�!�$��C��{i���(�ݎ-?��]�k�Gq�?�_�k$�|��^��'���+��3�1����"a�y%9lo��x�pS�X���e�6�'����� B���y��f�=�O�b��d�X҉7p����s�FM|1�����\��ާ3lbC�o��'(��t$�с��[O=N��*.��E�x�ě�����_ Q��A�66�L�Rd��^��g��k�տ8O�G/�A]�O���ު��-)�}�]���GC�QSM�(��8�Q��I��  �C����i����<��]�����˗�CR�N1})��8�{a�J젃n&�G�C��s��,���P��¼���xu�e]W.JM��X�ESCP�E{�"�w��VGRpB��m"��(�ϊ4bx��|1��E<��T^ҹ��0q͎@Y�_u�
<7�ѝ�1}�9�ɞ���n�z��/L�-�P������+؉�d�Q�$�-�K�DÒ?�=Fɂ��Y�h���e/�z�#��ܓ�w�
=kl�򬡏�n���lk)2qsŝ����lt�U/pz�3��(_A1_����I�A�[͔Un^�Q�T��y=�����W�ErZZF�Ð����"Ј'�(i�~���HI��[�I(UE�p�i��b(�z�p����d�;�@./|ԜC�q�D�{��%��2�{�W	�P�C���w�<�e��}&r��=^,��i�>݀���#��~:��y2!\sתڑ��\�Y5/ZGԹT�=� �����6G4:�ġ�m�/�o��~��p竖��Vɻ��u��i4��v]��2�<��̏����.�>�z��4��)��e��;~���>U�Z�CF4L�-\T�:}�	ZDE*���[3巢�KE��s��s�O׏r�v+����B����	����i;R�~w��)����a�/E	@�~�ҥX2~�}��8�"eү�hqs<a!&�]є�ߚ���[�wy�t_��s<�$�;��*c�CV�ٔ�lv�G��@��k%��^�xjZ�Ð�W�x�uKRh=�*�DN�����p��088��{-�2K@�j��u| �K�n�ή��1`��|/�g2w&D4�+�X�v�*w��:r��r����Lc	�R�חJH�b���\�C���gm�j�QJ���8_c���]W���Z�#���sMB�vj�]l�0�F�\w�]rI/�%�J�|@J��7��6��X�:}���E�T
�ik�eu/�$7P��X`���[ܼ��@G��\���g���p�}�z��?/4�juo�ft#ŵT"`!����t�i~a���e���	��Z���wS(@�ʕ,u;�������7'`��:��C�]���
��W?�薷Q�;�1�(��:.F���A��UE�V����p��V�ͨ�-\��z�ߗ��@ƃ�3��e���:�58F�`�#�m3�ߨ��b���򖹢YS�^��o'��e>�㠟���û�QWA��j����ɒ��]?j�}é��t����&�����L�*�/x?�O����'��/5� c4���9/V�-|��(N���Jxl�(�B��}���@!�/��xO�ƑK®����!�C�V� H�n�6�ȅ>� i�(��s����l�2^|��+�Ai�W�H-���I�J,Xc^|��{�N:����K�Y�[��T0)�M{��b#KY�5gg!�H��n8����b\�2����F?�� ����N�]#c�U�S��b��<=�ś)�J���4��D�h�ٗ�D��lD��6�ؐ 5���5I��ơKM���H�����>�w��[�t�)����$�>ǔ�W`��J��	�yՅU�fX�m* �=�G�gɠP�^|��M�M%�?���N�+e�Ti���d�O���[�S��'(T��5� �Un��u�n��ֳ��z.�
�p�L�7�50A���f�E��w�ůjv�"���O�r*���*��gZ[񆌛����_�G���P4�-ZƮ8�"���U_�.{�;��~?�+����uJ�8'ЦG���~g�>g��*,�����v��P	��`�+&�hl��>vFv�̐;H+��h��[���k�pG��)��$�����d-��<���L����a#�{�S�wp�d�D啽�Wn|�[��O�����`F��0%�G�6D9�Q�s\�ǌm��%b^�)@�u��X.��h�"�V�=f��( ���m�G��H+CS4�S���4/iQ�:��\N��M+��Ta��I�'�V�����Bu*�ȸ���!��!,����m(;�Yf���G����������,pSFB����}�;�㬻)�\���k#�g��MQ--Z��%��1x#��Zݏa0b�yC���v�u��kǴ�Y�j�� �����h�B�B#/ټ�6I�:;��Z�f�y�n����}B�Z��Q�?���ӽ�t���h��fm�5f�IYϳ��:L�z ���uG�T�Ke�mQf`f\-)�~U��#��߸8���5�*a
4��h��y��`x-�~�@����p�%��w�#�O1W��Sf��=s�� ���xX`^ N�ݮ���#�H����cms��b�{�f[����d�B �O]/7qW��m�0�x\�'X��'�]E~,���db��u��9�Е���N*9����h(J,D�t�^��{��a����b긆@UU��9�;�E�<f�h�*���:,�d&�}���&v|��~�^���_�#4n�?�4�_�}l=I�s�a���~�aű�%�B�#�A���c�W��ýO���~ �҃Z!���f�_$A5�f1��qC��^�vH�B&-9��}k�r�B:��w[姻��� N�.y}.��v�~ꊢ��O�(��m�#�E)j�N �0��]�W��Κ��N*���n1̓��<ja�����Ow�(q"��W]i��ռ��j��j��e�gyC!tA�N�hPP����j�r�,��$f��R�1iQ.���%5�SV���َ�s�,�L:�1��ʫ���d����Y��#�Ǣ) �� v�h�߄Mzc#�D����Rj�i2�\طd�x0�o�ڟm�"C���#�9�-�آ»����1P��f�'/֥�$�ѝ�b��;�s#�1i��M��6rjA���Oj=Q��i�����e�v<FzU��~N8Ʊ�Jg�5R�
�X��!�[�r��*���
p �;��ʗe�D�.X�А���]�J�F@?���'I�Fwi@ۘ���ǈ,���9*cї	g���2�>fm�j��=a�U�:�_x��H�nd��i���i�U&�a�ST��4�)���D�8����b�vY���#=�v��i��G����~�R�<o��yų<s_bx�C�؅7X�<y��;~y�-�`\ڽ2�ξ�<�A�[�б<ܒ��U�"H�n/�<HtdV�=���Ht+��Td1�����'��ڸ"�3�����쁁q��gD)����';f}_�xQ�ŊV�ą�F��3h���;vkXq�%>Go��8嚚��L�_�<��@"�=4��n��v̟y0J�$ٿFS��W-u(�e^����V�}��i)����eۄ����Z(^,���dŧ���$��Td�@���=P���L�~BrڅI��?���s�� �n�� ֏�q�F.u�� �N)��|�9��Wĝ寞e�-j�H�����}��̣�o*
%@�u�<p��ɱmM�gm(�c��â��	�"�4w�'�bm��P�c*�}ݺ#�?��|���?0gY���������ً��X�ϤVi#z8KI���b���R�)��Q�D-WQ����DJN�7�b�o���X��=񴁵�&E���/`"Cw~���;��w��.	`��ɜ�٪x���	~�V�f�@���1�<�ԍRFm[���p�<�X®�|E��(��|�d�fg�vn�IՆ���[�c���j��P�Y�V�����4�f�u�O^�����kV�X_m[$l��Wh�(�	a��(D����u���N )B�� �;����,M����`�
׶���eq�z��\����؜������^�m͎"��޹�F�)�u�K������9���6��*�lL���:���$�����톳x�S��� a(٧c�A�J���?}LA��ь�rp9���6��K@9nUiY�]k!�Ϡ�2T�zG��Z9n g��)ƽ`��*>�����}|��h� ��N�iWC�~_'���+�N\�WiǏk��>��q�K�Sv͢����`��²~2���ţ�(��,b���/#	�e��v��!~x��1�$5�+�S�	�H~�U���!��zF�!,*]N�K��v
��l��}CGt����U��[ޔK�&�Jo&��M����+��_0 �p�U� XZ,�i �Y���c*�p���^�QO�U����i�Ȁ���5_<���&��|���CVה����p�n)H�5W�R��Bci~�U֍�^��s?�gx����ئ���6��~d�ܒ&p�sq㐰b���SN�УB^.E�+�����ݚ���{�f�/�7/ �Q?I���4"5q��t9�봵yH�V�2��Tv�:�{xXM��)���(��dΈFp�B���Bؿ��怇L��6q���i�0鏦�=�0{ڽ7k�9�I>z��������I����A��t"���W�z�V�^
���~d������Pk���to�;��WQ�l��ap�Q_�.�?����1�2X������=�ͥK���'���GH:{XP�k^u��㗪�����.�K	4ʜ+�Y3���5��1�8
}�ߚ���rx	�����۞0�-���c�!��`� �=%��
X5����gC�������9�/U���q�Lu*)��uxv粑*����1p�´��ҵ��Z
�0s�
a����-H���:&�{K����!�E[W,�~AV��ce
����y�4���6,w�7�I�W�R���8^���/*�B��i���yC��;<d�;��[���>��r��a[w
�>�Ge�R����t�"y�j=�����1�ca�I��q'˟�V'�\�T���WE�fz�y�\x��DRc_�!���c�������c���5��u�/��f�6W���}�����~GzrO?5����~��z�����_f�c��]˻�<��`�\�޲^�V��h��=����4��ʽ�cX�ݩ��I�9�;s�Ԫ���lfE�;ڹ^^,U,����rf����ލW�)�
��,�9�,Fͥ�C�o����"s��_�I�WIwq0��?��"�?|;}��/�@��
b-��p�a]�����/-��M���nU����6f����U���ߦpJ���(��DZقS��p/�V^��X����z����qm7(��{�&��B*���%qaѐq��+� �(�~!�y,K�L��s������ʀ��M���m��-8����Wwi������,���KA9�C0Ĥ�*�q�J�d�$@��4�ٵ��$��ˣui�YZ,U������;T�� �!_D�WPz�?h��.$7Ӷ�q5�m{�$Օ~3�U�kΫK���Ǵ֑lf9`sm��\I��zu֑\`��P���3*�~3����V�+�e�*6=�@�R�a��\h"h0[�!��O���K�5�����~�D�A@���4�6m��I���nv =��霡}m�B��nR�*n�B�bˆ�����n_z��Kr���|3�*�Kel�}�M�f�饆.mF�O�H�3����/Rp��'\�����C�pr�s6�<T��K����ځz�=�܁O���k�f���,�˹%Ђbh3O
��t �^� @)'��Kv����e��>�Gb�HnV�II��1d��������u	�"��Z����c�>,(�hH����������^'���#g�꧎��>O���G��}l(�2��a�Y1��h�w�JpQ87�d֬('�#�=�vN�;�,=V��B=��5�f�-�)o��5{�o��w�vn>p����u��}�w�(1I���?�i<���< �.����hB�����
��lP4,�*�yVQf8�kv�󴋰]@��$�B����ӄ%9=_&S���3�@Ũ �q���) �4clkEm+2��Pm�͑CQr�i/���N�2���!fS�]6��<���ǌ���3�t(���-�&#�M;x��$_>]H�|T�3y�D�Z<7���5UC'ȗxs�;9���Q�������톎y.���5�ɢI����%��|#{�R2��(�T�N��s�O��9z:�7�>*06\�>YŎ/�	���&���S`�|�q���zHG�]�䔁{��t�d?�N���'rT�P�Os0�ڴ6�&#�ު� Xv $\���ļ�&���|��~��q��D��]��BU��У��}�/9�{u�|]���ʿ�v��8G�]{#�N_�ɜ��1Uoj�)�F}�N~3�l3�C��t5�2�#���
��i�/)1�^�T�`m�B&f(�[QB��9�l�]�l�ڰsK)ޫ���W5���"Y���k�B�?s������O
O'�V���¹�07��9�{+w���O�g��~�u�".ͨ��S<���]�
�dB�z��H)[�Q��T������B�̧M����%->�G�c���``�ɭ��f�O�1׼�f�=+<�%�|�(+ʕ�����rnµ́��z���k)m�-?=U���=nopI��QT�b �K7�.��ac�	�\y��X0S0�9����aB\(o_��_g���Kix�! j�q��}6g�x�V�2J�,xA�9cCA�B%1��i� �9-�M��?����GsЬXkqLD�[����m���0A��*o�/Z��N��D��*�<%o���j3y'��qy���>Y���7�O���
��jo��k�PK=zѦX���L�}З��uC����M%k|@�A�!�ʗɩp3������:�UPЪM�F��4'�52�q.����S�6Z\�xo�CDvȢ��g�U4�DUk�p��/YK+��$�{7�K�8w�w2}��i�8>Q�])(|N��A��HI0����;ұ���G�ב�#�>#TeG�`f��S ���盗Q"n��k�����]���^���/&6��$MDJ��Ƚ)��x��P�Щ�\ܤE�cr������en[e��SB@_O��L��� {.'�s�͚f��і.�H�OW�]T{Vô�h��'?�D^9/���c�2�Y�Tpp�	0W�D6�9泷�D-�s"�j)%`����"�)�S+�T�&h{V�_��8�&��w��4�rN���f�,�T~x	�2�"���d�Y��p7r�>�2��]'!��K�����$e��9��@�Ă��
�#7Ƅ�>���L	t�y�zu�m�y�?�J�a7��r�_�!�c�v!��C�c|S}���:V����&��C��8��"�}һ�ǵ[s
�J9��|��^���z,����)��2Ysoj[3j��]�C�}��%k<3�m2A���<�D*�!�M�(Qf�x���[g�n|��\f���{�:Z.X����,��f�x��-w-#�9r��l�mzA�o�C�x�#�����Z�+�5׻e��xl	2+1�#P�����%D2 ���+�������=kRX1V�/*mb�$�oZ���a�+.�WZ��ʬJ��P��a�XPM��U�9���� {V��zߕ��n.�]e�!ک�\<[LT݆�Yfw^��:��E�gR,���{D���ۍ��6�����y\��묷��qI�}x	�,�Y� �n�.|��e�����ӈ��@*�S�VODǙ�j3��p�?͓6� ��W���fM���s��	��|_)��[���5D�����&~hڔ;�WlA��m�Wx) �8l��3�GU��^#-|�r�)P
���ɹ���EOya0z����������g\Ӕ�,-7H�Y�� a.p����e�R��M?�c�qswOr�D.�̉馁m��s��1�8Ĩ�h��R�{+��^gY�#���<�%3�{}�dЃ3���c#�
tc���$��"ƪ��9([>L��c����s@���#7<�&�Zqp�4y>՚��Qa&��h�c��SN���d����B��X�絸�<L���`e#�i�r,:�X��ׇ����e�cyQ��`"���U��O�����/E({v�iR6N�fJic���U���e�ﬞ^��+�7�s��޷L�h)ڝ��9_���\�Gd��y�id=`��D&ʘ�Gߴ�+��@��� -޸Q�X+u�� �#m������l��3	��]������N ��Cfz��.2��Fއ�F�˕S$Vp�pqG�s�`7D��*y	`�ǅ$��=ƻ�U��ӱ��
�P}���*T~{v��$�������8k�D}Dx�hEֻ�O[|���Jpx;�`��l� ���-=�y��FrE�z�U�T��d}��ĳ��G���g�����b�Lc����Ⴤ�p6E�?[��\<?s����@�.p6ӛ�o��s�;C�Q�(�0�yX�Ym��I�.���:��{��ᢰ�9�Lw�yz�u��|_P/ Q	�q�Q����51��>G�P=�P�ۨG�̫�Ri
�˝���u�%��:�-I8��H��� >���+J����(���cƌĩ�Xjf<���>���HY���+B��P�&͞Xq�@���=.�:��,��;m��&�T��0q�jF�����!ؽ�E�C���* ��L8��.� ���� ��L©���,ɶ�ksǸ�/؜/Vn�E�6yIh�S#ql���K�e�<}��c���7��C;�z�]��ދY1�D�1叭�	[�O{Jy�����Of����1��4���`w�(��~�i�A�l�w{�>J��7|:�Ď�q�:*ޫc�K>ｯ�/&�)���[
���6��o�]�ˤ�4~B@/^��@�0�E����v�h���m�g	��� Z�$�&���c��wz{>H$%]����t��
���y)�>�}u1�dg�MMZa�C��J����SO |�2��o���ُ�����J����bD2�XL����^��@��@����
tQڢB$�q���둀�^�ُ�,X��f�C.�N�ԭƖktF6������A��]ų0���_���xO[5�-Z"Ⱥ`ۅ�	t8|B�q�-$l�W�,}�+]J��Z�㬨R�]z��~��`���Jv�_8.㢡����r�[\��7�����ޕ����L�5�>�o����5ֿ�2:탇����]�o%���7�A�O�d	`k����"Uc����S������!A\,�Y����mu�ą�R���o��.�͸e{\,lh�0n#��-����GL�� J ����þ�IF(� <)>t�`��a�
NL��U�6rw%��f��z�˿����qκ^Bt9ʾ��P�p	wAV$��(G.VLt��򅖆���C��M�o���Oml�(�����/뚕P1�Gf6ȵ��&�agj[�C���U���V@�`��s+���v"��K�Зl��m��:  &��?�� !j-�S�]N}e�r�\�ڒ
�������;v�F�`5 �r�2���7��X�GO�Ks�Ʊ%����A���4qJ�>��ɨz�bn�@��s�n�ν�I? ���F"��Y�NU�L���/W.���,~*O�x��uqv���!�PT�2o��Ȥ%gi+�]�5V�����L/�+;2���d�����)X_R�����.y2ֻ[�(#�B��pj�h���#,��W���m��G� ���v��v	�2�x�T��Mu� �-�h[�<��ȯ}-F�U��{�ƀK��b'�ܟ`�o�t?�)�5?,�-! �s��V��Ti�6�Hg���?ui$s@�`j��D������&!@��G%����E�6ܲ��>M|�� DҦp2��dȒkXj���
)������ -���N�����42�X�����c��V��z�&k5�s&�t�7�;L�f��p�4��ۭ��������Lb�Y7�fY���nl�F���d��j1`���l
S׆I���sw��,P�978T�?
�S�Ʀ����ъh��b	c��R2��C���H h`�;x����d��I�4�#��Y�E}��;~E�S��,�"{x��3�d�5UTXI��X?���dd�(	����t͈"%���{ZD)"�Jx�~G�S�W�8�E����lEJ`��7΢ A�=�d#���#VkN�8wF�B�����kw	��ֹXLy�ԉ8�O�#��n�
2��0�����И�B>���؞�A|�ĭH���[��l�r��=B-�����çt��d��Պg���AtZ��|��|�<�Un<[�Y����O5���%��rI�	�C�QC��r6�D�K����%uS���� K9̪&z��^p�]Ce H�e�߾) �S�������Ë�����֕���xD���#˒A��ht��(��r�V����|c�"�e&m�K����7��W:���͟Ἵ>X�����q]�L
��$��v*5�e�1>$f��IF��	��d��T:�����P��j��#}^{��G`�~����G�$Դ�l������`S��6?�kg�Zi��2z��8��K�Z�JɊۂB���y���N�h�̛az�N�g���) a�����/��Zq͏M�R�@i�V�h��K�O��w�Y�\�sh��>���\jjHX�B�*'�r�~�͏���c�Ƚ�L��j�G`2����r�'u� �86m'g4�����]��Pz�MU3��H<�,�U���(H!��2��M@K0�{���50�Vٛ_�n����X��}:ż�$+�P��P�䄢�o.O��s4�)S_�i� ��/���ɬ�ZG'Z��c`ʭ�K��t��GP6S���N$�*��?o��Uhp��n�ds�8�e�o|�����ӌ�'%wy̡`�'�q�5'ή1#N�B�q�˼1��5K���b��[�i�<�g�o8w��aY��:�
�g���ך0
:���ϐ�r�M���w�3SF}sW�t���]������}��'�~�sIFm=˨p@�?���i�����y�!b����C�k��Y]���C��p A&�e�%��78����y�v�&��-T+n�8�h^F��7-Q6}�,��lA4i�M�
�XzB��<��+b���}4}+�+5 ��n�͢۷��#�t羸|���BPL��7�噖�̡ȡ�6�$�]L�����8z��r�ǌ����!�Cl�a쿓}�z���F�Ш'���h���E��+Qe?�â���z��$����V��v)�C���9a� �6QD"���vm�ۍ�!�<ʒ5�[�ၢ��R
�W<Q��J�N�w#H���N�"�B<��
�	ƀ�f�.��m��Qg�9G�1���0�^�� ��i������ϛ���I\�ri;�o�%>�Sp �/����]+L���� ���7��҆�YC_fdx�=q��HK���r�/_D䚦��Ŝ�Z�	m�4tρ_bz���y|c�����W{sz>�F�{H7|�ܚ*6.��4�&[@�n&XŖr�Gɿ5B�)l��|���ߵ-,�P4�@��]i���//i�Mm�h�2[?�ED]}'����Q�v���Q����N���	�r�+����t;�y�-dx���cҸ�����׻(Y�10L�E������@�C"�P���Gn��B�F�r�����7$���fH$�֦��ޖ"����
/p�!Q?�v��Fq?ݽ�YAz /�	�8�Bܕ�Jio���Z�b[�D�aBP�{��@����}�C
c�_l�m41i��o���<uzr�k_�5�W��?<�dDNi��%�%���y"JS��ԉDo��y�{��!����r������W�̅�P�#����.�n�����'Hɫsc ��z�K��5�#Wz	*3�:t�%��<q�3��t3�cG�i�
�Jy�*q�"��y4#6N���m��_"x3D�d[�-�,j?�(�M`��3qb��Y��no���D��kjw�9	�Y4�sY�	����y�����("8-����g�%b̘�N��Kb�:����s���z>�up�m�uF�µ�5�i�%������|�~e�|Z�{X~+�aH��=�͍��1̋��-?nZT�9]ښ��Sbk �F�MtT��=��t�$UZoE��%<^���9����*.��n-i�J�f7�"�o��n8� �K/����k5��8�`�,����q���T[��l��4����zc����`m��?�Z{y�Y��

 ��$�ƌ�C=��"�,������L�����j�Ō/Cش���j���� �MG�$��ex�x���_@��~��7�`�4��0 {҃����W[m�L���(�ڴ�>�B��hڅ2�8��h�؏���f\V���MGV��1^���>�G�S���<��4����a5>0l^��U�Ň+W�g����`�7芅����>�vGN�Q�z�.�L-@�fv�Q���p6�@�r�F����$iH<��2*r� ��\��>��+�+ȍ��ra�|	҄C<�xS%U�!���3�nÉK���6mG��}�_��ZH�]/�uc��=�)�Eq�������3
dlZ�ϡ4���@A8_����i�#�vw�:SE��l�M���9}�M���8�Ǆt�����\T�ٗ�Jē�����ơ��5�>�5�'�d6Fʹg�s1b*����\�be�`����~~��1n��K���.; �xN'2�I�m�
�H?��]o�]2+�0q�P�P�j����46^O�K~Lg�J�̎0��]8S��bR7"eXy@�掻�HW��jD������?u�&C�[�r����oaT�ᄚk���
�I�a����(t��j�¬:G{�9 Jy�_�
��DӬ�@���*r�޳��������?2�..��Ed�P<�"d��-���<���6d�\�4���47���wG?o�E�Н�ˌ��}��'�o5�#,����:�ѳл~�V�"^���"���]�Ooy�� ��5�Y�"��'�N4=Fc2����e�C����X���$�)O�l	���p�Q��o4�2��%�"<픕ӡj�Z�����{c��)l�W���ڹ�$�W�����M%Z�2)c�|ק�����Rؘ�{��qwd�!����N�/��H�L$ҏY�m�V�@ٵd�Z'�x���=�Wa�)���A6D]����޿s�g��Юi��3����$? >t�\�,���XQĬ�b�~��~"G8z����aݸ��إWf�@mxEXl�nj����_{�K��@Lh�Γ^�d����W�mډ�6U���tfݥ��4����D�k��Jn�������U�r*���>Z�[��1>�@��K,�G��	�:��2Q�*0�wF+>��6���ORR��#,'_�H����Su��$�{���,K�g���6C�_'vď^��O�=�t"�@_���q'��CR���1ԃ�;X�1YG\���6�j�9�K�*����k�icv���H�ڟuQ��a(Rg~{���%�g:�N���@��F�5$>j;�����
�p�3;8�t���`z*���8����xػB]ۂZM�py��G��4��
f�zH5[7&����Ll��L����sY�H�U� �׵��a~�.f�O��>�&��N��n�4���⇀�OW#dk�At�0�z�;��Gs�ݐ}w�?d$wY��
_K��b�j��
�Zٔ�����������+0G4�X�tk�`�)f�֍��V"���D;�P��ſ~��%�Vb,���H���x��'(
M��(�Q���hp=�v&��Q�&��C�L�ƻ]��#G^����ճ3���Z��)��2N]ӅY;k�b����e��Ć �e�z��p�P�� � �Bf�_-�B�4�رd�^��'���[pCT�F���[�����ڷ!�Ji.V@
���a��e�㍆�1�|S뾅M偕x��8������͇��d��%{*tw{F
D�%Sa��+��V��%�"�R9����\��']����E�gj��"���4�F-A������Ehb*�w�R������q�V����\p�ܦ��C4���%�v��{;J��$�B�h�N���4�"}�κD-�w�˺�d����`"�CC���Jᢐ�>Y&�3P�Jz�n��� �X�s0=��q�p������L�����V�JR$1_<�����pE$p���zU�W�Xy�����B'�t�o\Z�]������c�f)��f��2�'}�P����=��f/��Ȕ��ծ�?�Ћ\rx�p����o�H�@��t,l����a�gk윙�����YF�cl H�����kFV�%�q:y������$�x	�T�fkA���$�|�t&�i���yo��2P䰶�SY<����~9��[�s�Ji�4�H���g^h�xձKX���=~	Lc�/�k:�\���h�k��o㍁D~eǪ���E�rJ���~��F��_����s�\�t H�A��ԡ�����]/L@�]a�kR�u�XJ�;yd��!2����D�Zpm {�����:"%\u+�p���f:�="�`�������`H��Zx�5q~��Q)U'����͌ H�+k�\*�a4m�QZ��qV����I���l�d>U��wU�dl��s��	O,t��K9�A¥:
���8��@~R�D�-��;��	���j������g���T+F�'��ʨ�fQm:n���fw��$���+Q&�T���I?<Pe����я}��r��𩿻�LY���,dP� �҅ݜ�������,:�B�\v�^��[C�A~7���3��'��N���H�7��+�R�F��l!ʸ'����� ��K�.����@�x�-�lS;'4X�2P$��eft�M{?V�i�y�#���"ܐ_�������k@{�@����AqOKRn
�28�驪g#L8bX�-Đ� ׵~�T�F�N�DM&���Rk��r&��`��9�S��E�:cV	B�"��f8��o뗾��M���%�����9J/-Vi7��=����`�����S}\����$�%�[��3���B��ۯOX���n��7�n�l��Ξ�S�`�V�yC#G�wz�c���RU�C���!wq��T����jw
��7~!+ͤ�9��84����>�5r%����%��-�r�kG㈰����	�]���W�>9q~��}�%C(&��VV��0�L��F��+C2�~տ���r������8�}L>��ᄅ�@�����Aa�&���h9u�*R<�8Vd,�{k�1�45�X$�������j8�U�y�Q
1��=`5ĐE���X��rn���!-�&<�<�۩J[=�ršr0�G���|�����̡oRa���e��*xXmkC��/�e���w��)�����]������Z�z�%.�H�
�͍
���M�#6�橻��b���ry�rh"@���f�ل�t�T�R;ḒIx.�h�"O�T����&��>+����I�c� g��^L��/�p���qK�9��x)��H���c�z�OӶ��)"��/�l�{������l��XLm�Dߥ����w>i��2�b��x5J�	�oy��R��,O�]�B�����3N2
3<[�U�x����Z��g�ꑹ��څ�!X9P0a�d�g�+*��i�k��eb���Z~��6~z��9��^,M[�S�K�#`���p���-�;�:㵧% ��BE|ZA����Sy�=b�b�n�o�D��bX��N��w[؜/9��=	})Q@�<3�k
7ËF�o�Aܨ�'(v� ��T�&,�P`>�&t����|���Z+ d9�q0����VL� ����6����^�n�����Ĝ�� ut`�Q<����`p�P?��9IBV�yp�7q�'*��xTɎY�l��: �tG��Sm�(md�R�Q��_�h�^v���F��I�<��:-��F�ʚ�4u:<��G��
��L+���B괻/1"��K8Ÿ�=Ԭd>K���$&�̥���^y�?��������O]�=t����u� O�,SO��?�c��0�Բ���9������gi��sh������F�a�I�x�ŋ�}Fw�4Μؿ+�#��yp�RoW���J�a�$��#��46c��b>D� ȶ'�S�T΍ŧ��m�����1N����[��Ͽfxz���2w$��.7B�{&������~�s���^����u�%�R	5�E�������ͩ��% Τ�7��E(���j¡!� s$Y�_�%�����O�h��[��:ײ]��Ouyy4��F�2t�r��D�?v���rՑӥ���/`U1�Yx�$���9�v�FQ��mFX5�$�|�9�
�5*�~\/��Y���
0>%�⥢�u�=ń���x�]Jxs�Uf�� ������&������n쮝���5E��-��grܿ�ʹ�\(�X8�ȈHhMF��^+Y�㗼*��%���[�Ҟ+����īq6�)Y�f�I�%��Nx�:H�Q�v����Hē{1#��^��f��zL���y�n�Q�A_j4��v�Jh�L�j��o�� �_W��FE���vl�8p$�ڶ�dwq6���XB8���/r ��p8#�`�u��Q�Ox�ݹ���"垩R�dc���8_2���X����)�,d�u��24
3_o%CJ�/�ꀈe�o��+e�/��I�%�<����R��sG,���Tَ�J�$��/������9Bh*�K�|�Zr�h �̑-"x�;{4�4���㝍��U����������mώ���y�Q$zj�#�n/��}�r��=��k+��@��>_+�F8���Wbk�-��I,D/��>�h����G�rJ���=x�`�iRz�CpBM~
�g�S�+�����7T�Ή��1��]?�<ܙ��%`�0��nK=v�A,��O�=�����F���|[̽�c���ji�y��ߣ�[s������[�jx�;�����#��"��,8�KC��SI[����
�+l6�O�������_7|�R;�[��'���e}#U��	��I�pF�?S��f�x�J�C[Z�9=涓�����y�=����d�N=Liy�\m���\��������(��d4J��$�^ƭ�Msq��`ȑ}�9Қ"���M�{�cl���D�
�H�ڦ�B�����gR'�% ��`�hs2�TJe��])�%����RU�������S�^N���q5x`j&�����9g�f�F�) ����n�>w!�G��t����8P6F\ڑ���uAH�=��Qz(�يh&{�`��i���z���I��/`|�*����-�Q�hJ
�e�m�m{��wA��^h6�(������[�*�2*%�Z0��*J�x�w>Z4z"_� ��w'1	 �^p�����w	��B�0Jl|P�z��{�	�&��+!����-���9��2��1��N����,���{UW�o���ci��f�L�����=_�QNl�C�+xHx�z��d�F�bV�22��g��0H6Od�>�9��cfU=q|��C�P'n��YT�n*�����������Uࠣ2���_v�x�Ǟ��&�����]N�E�(e�H�$~��4yQ��j�UTٱ�WJltDy�Y��e{��0�Rݧ�QVĘ��*u�bwI^�7�Z��٥:���g>=WoHtw�Ӎ�z��ُ��1os�s�q�%�K���!�?|`�.��.Y�O�A���s�2k)A�K���x�#��Й�(]�B
nXDS���q���?�X|���U�t��o!�rh�*���j�5ʭ�Y���`���h��=�+��;��v�'*J����>.ɨE=���q=o�F��.�%�2U�{ך��[��Ω����\�v^I�՗Ի!�zm/�	�}e{t�>Z
t�]���t��v�QA�B'R>���t����S5�Q���}��]7�)BR`���Mh_�q�A]��~rǞ�^��9�I7J���5��{�[Q��p�o�Q��>��l���2��Ge�d�j'6a��,a,ą� �n6̹%8ձ.]�?��1��ZA��K��F�~��lU�x�;�ꋥQk�c=��� ��SE�p�� �`����;
��P�qB��	84&c�K*�+�Ϯ-n���`d�:�޴VAN@���"�1�|J�i}���,(��a+L�Zy�Ӭ�Р�5����������+P9���1�Pj��p��po�<�ZnC��s5@t��.T�>.}]��SM����t��
����֝��r�j:�3��`T2���Ei�Z��n�4�>ҋ#��5Nsׇq_� y;B����}��&��M�������]'���� i'�QI[� �n.÷H����x,�������6	�� H�a��r$�ظT�,���+��\(������ߍGՀ1Q���q�w%��[���q(f�If�ėO���iי���+����uQ�v�t�P�o�G�^���Y�"���c������M+#�,A-��7�gM��1��5?2fI�*wD5�Q����)v�;�X22-�~���z@�a�������FRk������X(��H��8��������m�d�46����Sax��D������J�鱕K~'�(�8���d��2u���hh����z���>8����"ڡ�[�`�N�����6�ښ�(����e8��1��B���8��^���&�y�B�Ʋ1V��@�b�S&B�T�~���E�|�_�(*�����i� R��$��'i�}orO=:�4' y=�^	tP��?��$r�G�˧�l��I��^&�,cp����<~�>8J��r7a�J�&�ѻՐL��Pe�蹳�A���_k��^[�i]ڪ��(�_������_�X��ŤŦ�N{!���V���ƫ��3Ҟ%^ĥ
t���}X�9e8��ޑG���jo�ϰ��[5�K,��4;)L$��P��FTA��\*��U��y6��2͇�R����zQ�y��9�T�n�}|W~��e7�E�CH�.p���+RR��Y=�&5�l[����% �s�z?B|D���G�ۚ�uo����p�DC��kZ�����߱������
��(K5�+�
�ў��R�Wk������{$ }u�?��-�*���b]A�������_�189�%_���+c'5��x��*�P�hr��ZӤ�X&$&KA���P�`����δ)�T�jZ�\&eו��$�T<��L�%�Q-���#N�Xa�C�u�����sFv.t]>�%b�+3��y?T������򱦍�8�U(>����}w�SI�{X�'o ��r�`�G;ҝ�V����L=�%�m���S���)8i�LFr̼��邘��[:�a�+QH�p�a01":`^�hc�"07�I+2X,mf����Sj7GX�� ��\�"���T�rg��m�7;G1(��<p�$�זRo7o�|�d5v����ڎ���k� �%�3����	�������	i�W�
F݂G����#�-#����yN��i:�������&�R�U�#~ɨ���4��zX@��Ϧ��F\��;��'��#G`�"�t���!�o�PE_�' �}ɧ�����\5!�`�l2,`��k��v����]�˾�H���+��h�W{��4�z�^�އ��o��R���T?�B:4�;(�#��:�,�3��CE@Y�/#WIXv��� �ޱ���L�5�&Q��/�A(a����S���K���Bw�I������������G�]�Q�^�U_a4k�HA(p!�@O��;��0�����ZG�ֽ�I=�(x�H[�e{��>P��J<O�)����@��b�e ]�Z��@��|CO7�{˳+t��۷{��N)�ݸ�'l���d�E%���r�
�P��m��)w���k�x�Ã���!]��"�V��K~��f�n������~'�7�dS��q��"<Ub����P�=/{�$�Y��21��PM.�O���L�<S���
�~��8�0I���L$|��H�<CU�8% ,����4D[�á�Q��q�2������L#�gx�asC�Yr�6��A�t���X�,w0$ҕٳ`��F�"��^�u	��ݝΘr@m�Y'�:Y����c}ohO�r�דǏ�w���oo����ё_���%�Z��73Z)2�3��[�5��Lr���\X��y!���-{�������1
�X"~Vk45��P.I�������t��v���"��Q�
#��W��d���K�������]�L-`�dh�"
���EN�Im�輷@��T �MX�T���JGh�Y) ;V��吳����tﺺp%�Iw�sK4�Q"��C6�������jS�ㅌ�W(=|�`4��D(/4��ex>��L��4WN۶�>=�3$�5F�EG�!9p�2�X����5Z����q5�*���Ue�|�Iॣ�G[RJ״NƏ�M� �C�`H�6K��Q�;�_����V���2 ߅��]�Y�	��+��Ě$�,��i�6�� 3��O����/0Z��uFl-�ժ�!���>u�eE��2��
�t����ðV���3 �ՠL��� �G~�������0ouG>{�ȹPA�s!C,2rTh���� �ǎ���,�cv���� �K���
)dI*p�#��ިJb(�4��F�2��/F�W*����IjZ1�b���G���A�w�ۺ�h��WBc��g��80�w;
4>��#�便-�V�j�R��*���E�?���_c1j�H����ߝ&/i�aH�X��(.B���:��Dhn��v{ǞO���¯�h�}���Oz-W��/{!��~�!eľ'���P�́�2���DS�֛Rb{��&sn޽o��7n_����BX���@tG�p��F�=��Bk��܌;�~�l��o��9�D���O�ʹ�;[�
o��ѭq8lc�ƾ��Î���A~	K'�E�7d]�����>�D�3�)V"aw�F�#�~�<���:�b
^R	>�g!r;B&L0�����,���@��G�4�כĻ�-���wx�M@'��q�P	X��Z�DA�Q���2N2W9�&��w���i�l����Z&E�������B2��Ne�x�'�
��V%�~vd9J0B�j{K�^S���Ϋ�U�+�G���uɽ��Y�����=7�
z&�z���oP+[�X|�̀�{j��V�<�yo4�½~�h� =�Sc["�c����ɏ�|̑s8���P�.�TAz�>�"�Ec̲(�T���ޓ`�mC��9l��]��mf����t2��Yy�!
�*�|		LF$~Е�=��ͻC8mm���{9��u"�յ��h�D��Y��4��?]Z5zF��j�O�� <�E�S�:��5�$��d��V�yЯ6)��<r�l\˛׹:Oy�e�z����5�~:n!m��c��>�7�,Ɩ�6�M~pc
�PT����HE�Gzԕ��Ă<��4<�M��j���������m"s_��	�#_�!O�:��/]Q����v�Fɐ��i�D��ue</���n?�\_0��b�26���!�d�:�塟f��J�6�[%ԏ�^��߄"� *�L|U�V[2��]<�G���d�K�<
���f�D~���,>M!�@���!	��վx/��e NnN00x��Ͼ"e��%I@R�lQ���||-�6���Bs�%i�$ʘq8��sLr+�.@ǠfAy<�=�y���V�9�:B��J���)9Ҷ
��-:W�����A�	�-=x����}�%�x���
�.��.C�{�M�P��s��0����i?c-�0��$/����,RB�Ν<�9��g6�"�D���,��~��"�s_^ORW�� A�%QBG�vq���e�犻�
����I���U���֯U�b9�јX
�i�<�"|R?<6Qg��������7�
�*M�).@UC��\���t�`�9�}�c�\�m��j��w�KW�J��2����~c�R�bb>�W=F$[�ҰU�.I
��C��|�O�d\w(,ۉ����Omb0��lʝ}E���`P,ĵT���S��9OЌP�fN��{�B(�C��쐾���Xws���=�s���#;�O���62V���b0�K�71}�>zݥ*��D�9�f7����gH��5�(1E��nK�p�y��,I�� ����*4���-���!��s;4�w�u�]iw��Wz�eq�F��Ҥ���s���c������6����_�H�|�u)U[��i-/t~�L��`bx�*�{�F� h�V���{��� R�D�"Vh�Y>p6��M�t&�n�ˊ�����c��.�쌭 �)p_u�a�����"�U++���,�N����u�#�>��Ka��x����vڎv?{����=� ���Ed[+���M蝒@�C�����k��^n^�� Q��zfS�@9��F�]�&��2"��K��D�օy�G�0#ݖn	2�1\.0j�6�|���� H0k��U�TU�]k}��U1C�lnv���եҝ�G�X��_����o��t��Ŧ��jy�|>&@�©
�3����PH��պ͛��п4�����I����`-�0�Y�/#;0�e��b'�e�=��Y!�~7(�:��u<�5 ���+��
R[�A�,�"�90җd)`e����T�T��N2���H���Œ�L*���!@�VP���`�L��L{=ަА����Z��.�5�B�:���-bS�j�B%:��@��n�Hòq��J
r�7#$��Ŭ3F��<�b�����3�L"YC)g6��!{+e��%L�9��#���4MM��Tf��p�T��p5�������B�=^���)�P)���jXg�Ќ~)���4���Q�J�{���O�i>�}ݟ<�9���:)�ћ/E�^�c]^��xsLs��F�!���	\}�j�r\���o�G�@v��8[`Õ����Qv�xV��p���0���5l"�:��C���������9�t}��)��G�J8)��,FoLh�����6�W�~���JQ3��jVv:�_S '��/?mW٦C4�ܔ���sd�E�_"p3Y���'�	�Db_��i�6.)tr�M�nm�������@���@(4�N��=��_��)ޜ��a�|sU�R|j��_Z��[���Eǃ될P������"lAb�Pyꕰ`��@}�ٜ�������g���{r�s���"�:֢*�y�t��R\��tD��� {�w�(�'��@�x+Q�U����cr�w�Ė�g�œ�~�c��Y�g��i�����@N�mOO�Q�?7ۛ! Ϸ�I��m W
<�'5��6<�='k:��G�B!<ԝ^`6^�	[�=گ���I��:��V��K+�L����E-N��a���u�avZ�np`��� X�1�%ȊhQ=�P޵��e��V">؜���D���,�,��-�U���� ��\�8�F�ß��7�����'TO�
u��n~���~�-�l�� �.����L��ʧ`z=��n�Q���f�nAo��*qR��w�͛�<��ٖ�\�i���p�ɊP�D?=�[$���zpLEzU���q�����+&��zK�T���z�ѲP6SϿ2��{���X�b�I�X�X��"x'� �F��`��e2 W�a����{[�]�^X�8�TzU���1��_p���)lfc��*ђ]m?��|(�;�!5P������Z�d�����]�����W��!�u���n�?�Y8z��U\I�܁Y`βE"�;~�%9����Ǥ��֔=����m�Jm4�2�����-�����$$��d��Ǳ�"�	"/-U�ͽK�&2� �H�o�oqBx\�Swe$�Q1lhr"M!d#��[Ysw0rZۅn�
x�Q������r�0.}�g�,>8奏n24���0��L�[���C\w �Կ+,��<� ��H�zr?�;�Fd2{[�E���/�r]�ef�f��0�z/�^���<B�~�T�g�	e�֦æb���l>Oo�*�L� �0M%KE���@����^t�|0�����b��ule�'i9��<��/{
v��ˁj�Xf�dN�ԹD�jO�2��f�⛲�F?s��8�(���*a��L�{0�>���^�r%�v(�[�z���\=Ɏd��y
c�u�Ä�]�7`yc�mP���~�[֓�n��.�z��RO3B�z[I��nY�� :}P�R�H��? Gz<#L�K^�3��#*��ط��"c���PoWy�N�{���f���l�Ђ����""/;���a{>�b\ߙxX���H�T�m�ے
e�cev`�t�+N�B��}]��+�W˪�P�e@?i�etr�����q��X3�DN�#���E	O�-��$)R�����1G���݉�K�t��]p��3�:D�N�@t���?���-9l�Y�M;�D�¹�����:�_�H���6�\dk�N�G~��R|�H��l?ڌ�/�O߆'�C��O��q>[�ﮱSm��o��"F[�g��wP;�E;J�����'@�&�� )=���Y���|D���$ ����S������� ��zz� .2=S5���;�+���]�if���r6C���0F|"�,�L�/	#|Q�hfht�	�ź]�HK�u���=�P=Üf.�'�
1����o����O�A1�C_��ɺʅ.�i퉓�eqMh�����C�^�R��J-���,Bm���m�k�P���J=t
�2ɜ���z	�r��P�IK���L�d"+����e3�#�5� ����{�;�3���$��%�?x���� �U`��S�W$�����D�(�e����U�rE��@-�b�:��tJ������Z߶�v$c�s
����w�Y��!��Nփ����"p{��������&b�{^}� ���;HD��t�>�JF����&Yr�M���Ş�82JLj��4�n�z���ϖ�kk{�dǬ�X�{�(;���
�u@�$T	(0 �R��U����
X�6C�<i%���%��C�3n�x|��J����Dk������pp
%X����\]Yֵ�q�S��=���ẖ�ވl��h�H�c����L;�2i�����W���]��k�/��P��3���6�%��Tg8ԙ�Iz��螦$�����w��E���4��+�ݎx�~���6_�2qG�U)��SJH�s�Hu�f�nD�Aqqa�n[I�jrZ�ũ:��И�izH���g/��q_L���\5�*�ӥWW�g���s?��V�{�@y���^�1��Z�ևjo��r!"�CAU����x4O��s����k+�Yz���$�G)t��p��x��.Z�3ո�X&�Կ�#nsa�XL��њx�����6�E|ƨ^�[Q���hBxh�]�G���hb���<�A_mb@���n�C:rZ�?���*Zy\���^���'R�<�j���]�\*!nr���EvU��C:A�o����]3h�&	Q�;6/|�*1{dg9�Aw����}���D���亭x��M��(�)z�2�xF��b*��{%�>1,cOF�����E��1Z7S��������a12��Ƒ�N�B�!J���2���g��Tt󸰲�3'�O�u�^��&~�k�b�!n�-��c�2� K�%VP�?���P���P����8d[lw��?y0t!�@���KJn���*�ٚM��+}��:�9�Z�bت��p��R�#%z���^�q�1��eo4�� Br���`�賘oܘlQ]�lA!F�79���VۇzD�^d5����4�	ڧ9&i=�C8H"��=�m�� �b�Z��j:/D��wS�"��g��Z���Ǹ�F�ċ�S3!�C��R�(pʂީ>�[�d�����-�"����%�cZ�#,
��[o)c!����́K�o����9��?঎�g
�/Ծ����8S����=���XO���A�罽�]�Ex*��e&��ܛM��"���E�v�}&�q�,[f�Ҝm�|��)o������ޕ��3(���'�֐����O�*?�g���/i]ib�D�em>u
� �]�yq��i�2Y@��m+��%�_C�V!^��
�`B����p��A^S�5*�� ^�oQ�IS�Y�@�A��EB�}���кǊ�y��7<v���G�ë������������'��t���}o^�^���-�$�լ���z3�����r��{��1��P=|���1^�Wg�۲��ecɍ��L��&�Գ����``�eē����ܨ���*�G�ή�j����hQ*����	!�>b�n�3
��-�p�_�dýM��׮Q5)}�S�G?-#vVز`c_�mʱ���c�t1+���Z�I|��� DO>yj�V>�d#��� �R9=� ��cs����p���D����0��l�;��D���tlr���ֵd�"��鄏���>"�ū��m���Ԃ���J:��wb�����]Z�����Gb���G��h��YFO�Qa /�p�0�H�p;���t�xvG������ؓ덕xH�S9��f�����b/��h=�%q)å�7.Ƅg<�6��~�=��������fZm�<�Sܽ���La�/z����r}%��t,D�}���@�~����
��ٽ��&�O5��0{��ݗ��R�\+7���B�E�m� 	�@��w3ØD�[��U��yH?��C��ě������pG-�� g�gi�
m:_Þi\�	(3%���������<V�gدT�Zi^�;Ɓ����?ଁI�jy���{8��CXFΊh�]q1�y0�qT��������r�I��S+Uh7�fG�.��RHX0_�5�?��_�aW��@�,Y��z�8-�q��-)+d,x�/�[�	�	y���4}�4�X5��]���8���"/YRp-�A�$���a[_>:�hw5oH'��C�wzf��0�`x�������7�$�Ĵ�z�{*[��o���yW�Z�p���B��7�̙������ !��� D0���.�o)~� T�m�IX��5P@s̅�cnA�3���v��&��$}l�8���K��Gh�V$�����Bq��n�c�]_�{Q�i���h�������4�����M�!�dd��X���s�dz	��~��Y�@t���s��o�Y��P8s
L���6�ލ������Z^���A��������EӤ�o�~�>8~�;QoG5�[,�E� ��b#���'7o��RA��VSγ	h�G�ۓ@��S���{G"��`���h����%S'��#ae[D�^�ȳ9�C���h�����@ɛ��&a*�{����W�d��cݾD5�]Q��D�n������J3�F+�d*b��,Z7�xr�/�=�6Ԛ�;����]�����{�15��q,ʜ�ǉ��J�mĻ�'sB���fʊdrl��s(��l�k�\f�*��AM�7Je햛=EW�<�=�$���O@��5}cM����S�^Ű�1An�D����	H�!Z�s��eR�ឺo;s��N^��@R�ދU��[�/,O(��cm�sJW8���3YO��K��q/�����kV�
�Nx�ϫ��[�MX5�0=�:����uy���f�4wM .H����n's�&�}ɼϠLLM2��ۋ*��W&�ߺR+���=so&c��,���=xGL�$[�b	�ͺz�#�C>�:�$'��B�:oF!�+NS��X��s7M��@�������F�Q#m>�!�}b�K;kH���&�"��t,��|�E�6�m���4D��l�1Cj����.#,)ѭ�9Z�uV�vn��]MpL�q� ���
A�e#���<BQ��\Qe_Z2Ln�c���?�V��R�z��B]���}�T�I��q��a>&�,�"������^Nn���Y���(<���ǭ�l��}��_x��9Q�%ku))q��0��<�^u[��V@ņ�|�i���~K��Q�V�C�'���]��+k�ɫ��2�O�2J`��ZcM`�׌�`�ד͘7�m�*Uê����������y�;�̻�I��
$4���\���B�s!>'\U�1W�&q�F��Y��ݾ�d���92I���������o<1�C�(��s���.�a�P5i��w���d����A5(��d[(��4~ۋxcy׺���Q�djZ�$	 xR�ꈮ���aC���A�l}�C>Etfp�����U���L A�s2/׋׮��@��P^풿gc�O?I�.*p�m�^,��!=A,o{�R�u�b��½n����׵:f�v�S�A*'��_��q��ԉRC.��%lj×�Q֊�|��,M�㛈�z	��oMXwa%���l�ʵ>�h�NlQ4l�������xbaerG��u8��)l���_^ ����d'�&ݗ�	�G��VPzOdGK�V\_c�������� I�	��!�r�Y¤07fd.�r����k��6���X�['adw� �X�)!h�}R�w�g�����1=��O�e"@K�7��8�uL	
�d�&�_��;`�R��eR�WV u�\���X�y[�oe4U8ű�ܳQ!��?�ʖ��j����W�~?�N�ר�����d\���)���v��MA<��\9Zwg��&�8���έk�����u�[�!h��C�W�H���k �"�<�4ݱ�\z����:Ue�3g�s5�ϣ����#8_3{����.�]�W�d�1@�������([~L�tB���[1I.G��i*�6��I��p�j�a�p���:��cBe&e�c�V[.^ņ��
{����&��h|���c�S�q�;B��YR?|ȝ7	����<�{#������������T�zGכ{|���d�m{��7�wO	^�Q
j��=#	آ,rK�b�[Ǣ��96HK~�Z�N��0Z�60A�F�VC|��dشӇ{f3Y����C�����8�#�����"�TeUJ��F3�.)ƣYaW�ƈV�1Q��f�,�0�X(GRx{�� ����߃��̈́�,W��>6���4�r�[9��*�N�~)޾�c?ZqAXI�|���iT���/g n�rv����a�i�>�!c�"������x���F?�qQA~��Xb/	��a5�Z(lƝA$vҍ���d��g���&߼6�~RbJ	�a�WN}ӑM����rq�^6��ς�ߝ�çO�8���=3a��WU���m;Ŵݔ{��y��q�� F�nv�}pQi���.͂��s@���p�Z�����~�
�s����I��r���
��|uHx�O�5�X�+r<�޿@��ad���U*�����,n���Ҿ�\N�;�[i��g%R�������R��@�����
��;�JK�]���0�t��?�b�����F����Æb0�_�%h9	�S�5���H9�m�'�������N疠����9�av���L�̏���
�����9�՘�И �����I�������2�p�
�v���񡫗O��r���̊�կOO�* o����pP�d�i��G�G���9?��9���r|Xp���s:Ip5�5jݗ�/�\���VƨQ��`9�y�O������������x{�I����(��(��`:�ҧ��:lo���x�1�ʢ�����)7�R�c��j�β�=r����4m��Z���$ ��x_��b�����<�Eѣ�.��}�qI�!�2mzX���]9B{%u:7�{2�s��3�����c�I��K}���I���$�rI1'%Ϟ��}ˮN�P��� ��O�y�l�'HY��M��Yr��"]�q# fv�:�O f��qύ��g�䲂���8�J�xo�i���>�LV��?��:\����"+@���E�y����b���B�X0J��HJNne�;2�" kzL�N��t�ٸ��ƈ,wK�CG݅����D��$]3���''¬��θ!TK���m؄���~�j2��ɥ6DG� �!w;X4R���i٢��݌�Z��
��|q nԨ�U�O�����M��������AZT ������GD�pj�=8Y	�}]�Mݵy5�$����*uz��6���fyD�u���5�&7�n�y�B�9���y��Q����Qs���Û�]�6��t��N�|	8���U81��nD&�"�jA��A�H��+�+%����!>)��N'n��JO�ɩw
u���K�V��p�H\c)JWU���DvA�Ȳk��w��ǐ�b��c���G6M����.��,w�.�$�P�rU���C5<������Q躹�,ZGuC����%�uG?�99� *�f����%��
Š�Pɏ$X�gRkރ6y��������������n��i�z�$p�w|�~�W���c{��>Ď�̥	�~PY����e�^�6l����ҶV �"vs49�#b�Ph��]�p���[u�=j�@���mP�ꩽ��4=����h�6���$�A�pTrjw�n����d�����c�G�٨ `,�ˎ&��������.��A��(=)�}h�K�"��Tp��C
"֎�L{�֡q�\����w��gD����w�
d=3;�+.��`<�R����zL�"Ǹ�
�x��������*/�4c8o�w1$��Z��lm���g�^����>
a{@�3���p�V��ڬ�?�D�wJ�i.i��0������3txG���D�����p�e �{��w��D� @�1��'z�3�d��jL��P�u�M&��M��(��+�;ʑZcZh�xb`��9�JԞ�u���.:3�W�G�%�AYhs�,�"�ɦ��Gi��*���@:p5 ��z0LX�Fz�����d��<[L��hy6(�S���" �ш8~�g�mTE�݀L�y�C�*.9V�a��&=Z���hU"�ʓ1�v�m��%}���;�/Yo�s���qZG�v\ʨ���`A�����Д���i�-��=t>-'sUS��q;k�V�q�J��:>h��y,���uc�W>���������f�(�?؎Ɛ0�����Nl8P�ع��%����c�w�3d&[X_QWr �����4����%��{BRǴ2�Z^�}n�Q�>aW�����G`N�H:٩�ކ�l�䩑�(��yRP��)9A�`s�&0�%�.L��e�� '�7 �a���a��4$:<�a�����C-���tLdIH�k���A꡸�� � &[T�����V	�GCIݬGP��sO��D�� ��f[�bۍ3�Ǔ������H�x�T�j*?Ճ�G{��p��˃�]�b^O8DN����i�|���HQ����~q-����ӸÒϽ)�B�]
Y�8�況pk^��� a���7�"��\9�(�1D+멙���K\�1��6펮�F���kq6��)�|�����b^{�[�=�K"����-%&.R�XsZ�T$�mI,Y�<�Q�m}=��w�X����1Ec�;���S��;Id��I��#����g�N��GG�R��Т����Y�� ���p(��M�������G�Y���������h�5�js��I|f��>T�!w���.�ӢJ��@w�9`&PÁ4R�K��>�ᶊ焸���'Q�!Ż���^��g� ��u)�`1����6�0@�p��	�甴p4w<�ycPj�&���ח5�Fш�l��8"i�O��0[?�ɨD����M_(wM�ҮN;���:��)�%�f�tZ\8������\��x�q�U2�RJn��v�<[���/��w�~�P8�v0��.��i�D;����4Q��@�*������O/��r#�.�r1ˌ��@���������A3d�x^j"#u7���iKIT��R����g`%.G��VY9�AC�jc���`}�F�q�AUӬ<�(���"f�ƏX�6��vQ�<;�n�c#Yp�j��[�P�o�;Դ��	���E�����~�yn��l�Kz.�8U�;C�Ӟ���a�ioɥM��Ɗ��V����3y�Ӑ0�.�K���߿��ꉆ�b���w1�v���+������H\A
��:r�c��H�qP��_v}��CtG���3��t�b�s�ڷ���l�H��j��OZzFBGҺ>��R�1``0��U7Z������#�4��q00oÝ�A6amT�`��X�_�qw���F@��G�эIN�2����fy�R��>oŁ��U��[�ӘU���B˹��E,���-�Y37���t�������Oy�#ҋ�Su)��i��'s69�q�|����Hy%c;L Vf�E��;�c�}���ֆ��bq�GP�;l�ؗ���s�oO�\t�e�kH:����\��Ag�S���ݜt�Gdlϫc���������u�@��99 A�Sf�6{'�)����˘���Uk��n�����M��cY߶?�0w�n�41�� ��l8�;�ڧ��܁���h����T���`���u	�NubHİ\<O��4��i[е]�`�:����a�s�O�۳��3�ǁ�p�(����+���(a���X�6K�-�x�xg��� -e\�c&�{�b�߄́�����=�bl��
,����R��⎼3Ae�/�7��Ru���q#�\؄���4����7_�O������]�\���P1����������\�r�F]]�"�E,/��=��;{��ґ,c4h�cj���	�#���M��E*��'O��5�h��z|�{�6����Qg�'�.���3T��4��+v�se�c~���*����j:��`�h�=
��B|�r���W���iGO0Q]cƏ��R=%�u�M~�fg̻*L��<���qJi]��� ��g���6� ˲n���FG�[\n}ћ��Y�-���D`�TH��Ka��7O�e��+�?-
�h29q��1�� �1����&F�l;�^X�
�c\D���	���<6C1��<�ri��EP^Bt�k�2{�KOc�z�ŧ�m 6vS�j�.�9(����c��%Ɣ8d��Y~�q�X�)�1]���`&��\�{�=Rq#6��/�+�!��/򞱃L�#�I��JTM�vh	�R��к{�[��7V��?-L�2N�$�uQ��m��q���l+'%��~�C�+�#�`�D��Lm���"��*t�{��em��@��։j��c I���edtz������pqiU/�I��B�>Z%Cѯu���b��H�Q4�5Cv	`@*�z��^%�@�xT�kfv�٤<W���!��b�h��L%��Ŋ�yc�r�K}�=�}��^t��'1�ۜ<����9��p�6�.�d��Z�l�gS�r�X�eF.�Ü�}4w��&c*MD#�PC	�`Hj�B͔�CW&�=������^��z��(���__�.p�q^��O~����8���Yc�N:F��ۭ�0�X�պ[�X��6.7	B�g����!}U*W�#~k�2�5��l�y�|��l��sX&jKluBCF���{̑#w��Mw��6�1gL���T]���[r����o����Hx
fM��voiV�|N2:#�����s�UAҌ(_ܗ34G���6r%��>����]�6�\��N�~�'�HcY���Y`�D�ԵQ��\\8��P=QӦi�/gl�R�%6Q�Ps�2f��C��C�GG(d���e3����j�}mo���oD�1��u'�/��,��M�b�yQ>|�I®��j�)���i ��~����n�ws��%�WZg^_n�\�z�kp ��1E��׳���`y^����uKg''R��Sv��(�g
��{I���bAU�nԀ
���Y�cmtE��o�������:P�bW#�B�V�+ml�=k�uC�_����AaRk�ԩ.���t�YYV�p�I��8~j@,a�A�C���qf��Vi�̱/��x��~����"��uu*���ϼ#b�PH��D8���3J�.��ա�<��0��p�s�e�ж|�f���6B'�o"rB����I#:K���ߺnV�[�c{���`?�����^!��k�7]�VL�Fn�I���XO�W� �F���7���ǝ�f���/f���H1*�$=�>X>:��B-�Xf0��~PҫŔ)��M�_��z�~ (�:q�q(�
���7ݬ��uZ����(�'�?]2V�߿z\��Y8�(��Z�r��a��8^�=�-�Fmņ>In|W�yF���<�3)�S%~�P�3(1G2W��'5}�l��#$��rv,(aB��JZ^T
Վ��L�� B�ϫ�y��h�x���2�K*�*��b�y�W%(
�+�^Ju*����)�����rs�]����mz��9M.A!@��������'E�ɪ攩(xK�z�߭
�"b�P��vS�*8{�+�w�zTd�ת��������u�uWBT��}dxE{���|"�ׇ!��V����$5ڭEBnk�N�zTr �Ă�N�}������@9��;�l��7�A�p��U����"ޡ団ν��[tu��k��6K�`ױ0��-'o��\Crp����"���Z�^�D�<S�@�Q}�J9�J�͏�0�4�Z���:[F����O	y꩹�{�b��P⣀2um_��!�yMd܁cFf�oUK�]��(;w����6Լ�ӅB혺H����~R�3�B���;����Nx�l��o�-�O�BHCu��r��<N��a�DF���r�*��2��j�%sη�t�~(�n����-�j��-ʉo�܃��OSH�W�C���`��,1��c��H��(�ܮ�z��k0(��p�F"�pB3E����$]$�����ɱY�ᕧ"2HMب�jk���4�V�mxYi�~�}I�2�Po�[������ʞ�+v�:�Eo���j	�B��Y劶������Q������0�=�)a<c.�(�Y��C���T�D۴���ߞ>�[1���f.�v����)�][N?��5P���6>P���8~��ó���I%���PJq˔�E"qz+-J�ol
����n��vH�R�4�:L�q��2�1i�|�BL�ye��`����Z<|�3�e�U����W%�opQl�90�A��~�4S�Sޠ,yןl�`��*�5I;���*�?u�����_e�_C�U����i�\�n&&u
c�C(F\�aK���!���)���?��t�C7���ȧO����6�0q���$��UO��H>��
`���Dǌ�
�c�4&�`Q����]��p9��L]-X�N���W���F���>����R�x��
ǧ���"W��Y��a����ԩ{��kB��݉C@�������@�/�
l
��ڢ���������d�v��ON��09�Z�AX����m��1k���&oj�uD�ԍ��-��^�~��:p/S?�N���+*�J4n�)���P��J<���9���^NQ�����b�[6��"��� Ow� ����ɶ���L_d�C�\�'v�,f�E]�RV3�R1���Q-���:�!�.a�IB��8�S���Vlr����_��L(���u��6QE�A�u�Jr9M�n���c��n�C����Z(�E�L��gtFEfN�h('��=��BV���v|�=�	�������t�1h۞hҸ&�L�[���A�4*p�>:J�x-o�2�	@�WK�Λ��Ǡ���7!�*U���*�Zn��<��ҟ&0���7>��0�(�M�	)�`����|���������&sebY�2p�����qć�2��Ql�|֘�vŒY{h8A�r�#mg4�R�ꢾ�3�1�	�$(5j<"�]�~Ǒ�p�b���nk���\o�]F�ư�z� �����^�Z���@c�������$��N[:���l͡uz�6��m�.����{zz���)��3���UHsfMw�A��[����dj�,��7K2䴗�2���J]��=I�F!��]������K�E�sO(2�����k�����(r�dV���ڠ�	�z���a/jqy�
�M1
z�%F���mt���I4��m�O�̘���C��K���wc�/(���5��&0��r����ע�$ddv[RZ�8��5�x����4��k��rx�IZx���r�,�n�B��� �`H��@E�$��pn�}I�_K룹����u���-�	�>�v����ZZ��������(Z�(�W��h�9@\u�?��X�5�`���㞐Ң�s�l��H},����"�݁G_�u` ��nݼ�D���D L�9Ѐi��qlw����T�K8�tAM��HZ��&�.s����Eoa���
��6��w>�؞�h#��n�$E�o�ѶZ�Ǌ���:��N�D�T��oN��>fU��h$��S�m�e������ޯ.�1s�~2%e���ͥߗE�'�a�|Z+�5̤L�1�J1���Δ�S��R5*II��v=�ϲ�G�+�8�z��;l������DyP��k��l'V�yו�<�[�����.N�+G$r&��PC��%2d�5%�
��e���QB?�ڮuߘE/�m�L<��Ӗ��J�J�Ԝ��K��!���pQDi�p2����F�Y�Պ������m�w��������+ۘ���	��Uzb����#^ux֏`��K���"?ž^l)챗�-N���W)�+SՊ��]8��w�Ei��`_���c��>��e&W{��[#S2��T�x�1�n�kbYv��VΪ4J�B���8g؁�Q�ze��.\��~I
�m��$��}cW�D��j_}�UFF������}�%�\��z"	���I
Οs|;;�7�b�
�ҪA6�����[vg:��a�r�:��PN�m*]l{
�^l	*��_m�gh�l���W������"�>��	Q�7ǰ_���?��nqN����2��rh#U5&T
�}�d�}��%*� `�����5�O(�.J._l����Ƥu����`M�hd�łZ�`g�ߝb8ъ��u� ���=��c_�H�0�i��H^h�8A��"���p��Y���F�j�PBI�w�8oF�, ��^<����}A[�e�0��qߎl#��-�.��s�Cz�����Fw�pɑ��÷ƥ�����X'�D�2��@�������x��.@Q�µC=��H�Nc�%߮�;���:�<���`��O��W�m���08��֠vV��*��0�d�d��7\n꧶][ˢ`+�ACVF�S�e�����4Vf���o����[�,�������L�4"ѼB���/�@W�v�5&��K���r�������\8�G��O+2�q�uM�n��I���ᕁ�=�ا�(�hO��T�N���h�`3����24K��D:���4��f
�����5���hk��,�O��S���=��y-�\뫋ث�my�OU\r!��>�R0RRs[*yŧx��:����:$/�	Ҥ�b�hT��B���J�@"Z�6���h��!�����s�oi5���4���.�mm%\�<Z���&�����2M	��7�)�H����������ke�~�nmp)������ュT7�.�0�l��n�$��6��9���b9c� ��ݛ�]�����`r&�β�7F~�Z��:�k'��7FZK���ܖ�ҋ^\�\�Ƞ4PL�����Me��@�r��@���z�Tb�خy�G�v����ێ	��dK����.K��P�{�X�'~F�O�D���ϭ�RJ��Z=�hH�#��B�m��ƭ`�ү��G��r�JK��>���c�������L���'�
*1�p�F[3�S�=Zz�:���	Nݿ�34f����#����@pq��Nn̼t.:8��;�����/��
��T��ʳ¿޺�%`zE�'ӹFJ�0��YӍ�熛������K�\�
ҥ!ʍ��2K���7i!!9����Qٜ�ۉ�`R�Z��et��-�P���1�&@�����c�鄞ɬY��A�#�eC��\�p��t[�)��xZ�y�YM/�]��'�V���R|�� �-^Mм�P+HL��+���*�����X�u�t�^�ͱ��B��o�eU��K�jp+g���	������FOȍ�t��W3�԰S3�b?]��q���1�	6�k������<�`	�h��Q����+$X+��H�1g��P4q�������Ph�0t�Ar�լ���5I��9�Lt0����u&�m
M�1�]$���r��+_~*F�X���+0h4ж9� VEC�@������>����C��,̈́�
����^����N�\�t<�3���:��,�]���i����|� !:�+���{��KOϸi���rv�����C����������=��Qܿ����Z4�ZHCz/��%�Y�����`k�Z^�x؜X�6S{��=��ߗ)aL���ޏ�~{}����uT�T#�����'ҧ�rF#Z̭��@�����'C Q�[�a{�����K���b,Jf�6��7��;3�v8#mdt�i���[��.[�8҆X[�0�����1�Pq�Fk��ݯ��0��TLP�v�@�K��C�E�xq���;�[�FB;�"t>����vꙒ��Y�d/��ZN?��B͍�.��	9��������څ�+!ym���F�3�5�E��ߙ9��cB.���^<��Vg@ܑ@+Zb(#�,�Դ(ȫL��'�[jU���*��4n����U���#$��� ���&���/��UA`;�86��tv���ᘕ�����qK�Mk�sR���_��P$�n��)�eN��kD 'ې��i��!l��D
�X���V���4|��m'X�_�3���ϐK��w��^�s"� "w*-���%!���Y����}������'��B���s��"�"8(��s;���/K
��e�q3 UWEU�=���=O'a|�t '�8R���k#|�g_��7p��� ��#�.�#���r��?�Cu��ϋ��"�Nb�:���P}V�3��-��n���F":�/zkY�3u1p)�l��[���IS-,���{Ӱ��B����bףA����xS
�Z�ݏ�hrX]��y.���U�v̳�pϑim�����ib͹@Z�,R���n �@���1Z�a��f	��!�\#���Հ�ۉٵ2���DM�S�.�٩�Z�t�`��j�1�])��Ǐ�%��H+&��	D�@�dc���~1�H��u2���l|�VU��!3�"d:GB�i��Dѓ�Hs�+���#�u��L���`��xY��� ���K Io�U�L�࡙��L�drR�c����iQ�=!FFߋ9�3�,Zj��ƜT���!JQ<C�Q��߫gе��xbhw��È䜟Ѿ\�_L؆)̀K���l�#�Y)���n@"#�:�2�ێj����
hg���d"S�qw��{:��:V�P�D}\�X��+���{����D�|bn���4�ݍ����Ւ�u�(dm�Q������?t�i���Psʙ�7���pL���Nv�d�p�:	>�N0��2m>�U���M�TXb��'0�ᨗoJC�#"�g.���u���PC�zo}d�b���j+p2X�U��.�3�פ�$��LKc�����DM�Wax�8��o�ʅ񥅘�쿝g���%o�h���� ��2S�iT�A������R�A�����)V;Y&|�vi413U�m���/hI��PՐ
�T��^�y ��e�Ĺ��81�}���C:���O��-�F
��
�'����&�jf�{���$�-�r���G�`;����{E�39�)g��٧��x$���:"�~��eaW�2_r���b+��r��(���F�u"A�Zd�{�$�}��d�Tkj�7�-��[��h,�5�E��]q�zz4��yB�M����b�?�p�O,:"B�F���� [��`kvQv�p��Ew+���e��_��>
%�*S��7�<r�Y6�열z���$��Ҵjr��X��$�Жc�V��[E���X�'��׆���Qb�ѣ���G�����]�B��(�Q6�<^���'+1�q�S�vl���?Mh�ZXd��a���"�|;ϲ3��®�;jL@S�@�5�e�3��,�^o,,���	uIU��n�~�d�y�rō����I�)Χ��ֺ�zK%a����m��I��=|&��#�	 c��+U[�4=�'/	7U�كf��T�Z
�)��*L�������4zK��.�X_��
�()�IEX����k4c��g_��m�	cMf��H;����5��7վd�V�4�_�H2`"hLv, |q/{�ݲyi���	ΰ_g�I:͛q�� v��_D�7������3AL>�53%*>43?Gz<Al\��|D����(����t�Hg�w��"��ʇ�S���c�1C>�Q7�;����&
���L�!ʵV�GN�kY����%S���y��_Ra:}�>�;�e�qW�藼st���$s� M@&UÜg_;S�X.��{���g�?~������AU���8�-ݜ0�Uo����N�y���cD��vG��<<������!B�m̶��;^��i{�R�s����iT��زV&�&y9�E���fbc}<�.�_��-�U3��xmO�;Ɋ����V�G�g5sA���6��Q/��k���}S�G��hM�Y/z[�t���FQڤ\f�IPX��y��"5\��o��ͣ �����V��s�P3�XfX��z�V/,��+O�>��ҪL���~�敉S�8��H�py	E�aO�To�ڕ����!7�a�H,�� �:�\m�(�F��$ê�y�,ďՃ��|趒�#����Q�U�.ʍ�&�p��~qL��;�Ǌ$��ɮ��,|�$0�٭F�~�Q�HΤ����l6�r��50�3oI!�\XO��!����T_�Xέ������ոn��\�f�[�	�$ۻ1��.��Gg������֓��Ubt�X�ŏB���@����E�`g�CC��>�����;�,^��FM[i�X]�/ �EY�%:�����l�ܜ��ؓ� �4Ot'K�ۮx��c�}N}�E>��5����' ���̜�:h�&�W�����m�áe��e	̞�yVָ�
8ʙ��Sv|�q��ʂ�\q�{T�yb����7Qj���ܤ��5�QE�	K4+\V�2�ɾJ1rD����y���q@������U�2	���Ҷ�[\���h�4�sڱ��`�PCfl�G9��lր"����孇hN�\�![ش}I�q|,ѧN}F��rOy$v�X�M��T���q�N_*w��vi�����I��t`������Wއ����7,m��AKFh�ZS���kR
��M��}�FfD��zփ�U�� y[5�}{⃕fru2O\�ӱ��j#͏��ZH���y���+��٘؂�I�k�Ƌ�@F>����^�A�I��Aꍾ�3�8�@����;Թ�=4&r����}�^��Sp&�T�����fNV7�z��W�:<}��Q��LiS�N��:����f��魶��ߨ}��$������F��F!�
���	C4c��d���}F��T�O��W�2"+>�*3@l ����%d��h�ӹ��hBQ �8#h�[�mr�����фk��l	�:�+�>m~Q�87�\5bk^�
|�� �b�a���qq�6�Qú����T8��<	D��9<ƶj�:��w>�*O��Id�=�y~$��[v��
Kc~\���Lr.z3B��9OO��L��m��`��\��,�{+j��ӌE<pł�x���xHwʟ��&D���3v������`9Đ~"�s��h:5�8\��8mw�ӳ�}6�C�֞����%���Gtt�j�+�ӌ���q�k�놏�:ce��: ���c�!�J�Į��� �6�'�r��BS�|�'AXX�{?p\��n
V^5"b2p��f��o�i��۾)u��Gԗ4�	���t�M-z
�+����Lr!PZ���
�:���d^��|��'�߄������6�#�kk��B<��?�7����FH�p��X/�l�DK�qN��M_�.�o&���iS ��a�j��ץ��9U��֢���9���%xj�?��eI-m}���#�`"���T!��#6Y�Ǚ�����n�d-��&1yD�hVjw|�L��hWBOM,���jL���u���r�r��eg����Wt�qS����fGo��-�aJQi}:�$�F{�Qi0I�M� ���I��<���g��sf�ߠ���7���0�U�X3�\��4/ʩ�$3Ĩ���'cb�ѽ�KU�}.b��W������� z��6�d)�H����Vrfu���X1����- �݄���R0�5R=�.qf�\��N�g�3�wxq�&�GbHo�sk=c��|���,�HJ��B@?̐J[�"�G�CܑV�	.�4�:�2��M��;s��O��V~��0��w%�?r��	O}��`%w��|��H4M_��������;����dK���r�JH��������'���+����O�Ѧ���J���w	�Kt�p����P����U����dh���f� F�b+�X���Sx��̘�-��-[Q�hҝz�%j�
_YNѷ�z���#���UQΔ�8�&j!]>l��+�(ך[�j��1��<����س���l�;lM�m���e1�Ĉ֠'d����?�L�G�X����r�h<$'�q���=+.��L�"X��B�� ������3�q��9�N=�GX^�v�N�X���.��m2t���N(d�m�e�ـE��\%Ҋ��b���8�.FEL�y��?�,&��L3y 3��k���� #���Š��½��Q�L8�h�82�v�D?!�dmS�	{����
��G���Phޟa|�Ag���GXHc Gpѵ��9Sp؍~j�%
��M;,5�vm5xI��PJZl]���%eM~�n �u%i5I6����C?��T^Y3�E��Hb��C��yl4� S'��r���(����)gi.�_�ռ��/�� ���5�[�Dy�;���b��a*c�y���8�xW���N-4��������;��}8o����0�7.Rxbq�(!98�u�&��0�16�#W�4Y!V��?�/����s5��vk�ƍ^{bА
��G��C�=^X�+v�J�1����g��j�(��(x�lɖ,t��`��Dk����i+�BjH�3����W5�Q�]��T��[3�%�3�X�����2��4z��P+h�c�ɗ�D�G8�q�zK�|�6�e�����q1��+w�ؤ��������ճ5��+>*У��Y֗̈́L$Zt���oY�q�E><����s�ؙ�jv�"�nu��<Z�k��@&:��B���̟�29M��^�W����{�{kVY���O/�� ���Bd]�y�I7'��#�J��)w��/	�ր醯^�N,��C<%0�D�
�Ư���7#�	@f����c[��
I�36�ά&Z�t�<�d���xY��I/��5֞�H�{��J'��Fͼ�3�����E�.5�P��Xj7u���X�b�	�2y]K��;I�i�:38����y>5>����Q���K�T�`\?Ŵ�ӡǳ����L��5 �%c6j4��h�yV?̉h�����:"Ͼ��N�������)g |���ǽf��{�7d���h��_Xت�@|�E�xz$X��4�iu�����_�(w�s�R��P���tm= J85b�huw�Z�p.Y��a�6 ��qh�Kiny�#�b;�o2Uw��
n��!I}kR�I���p �+;��c�gq��VUV����xx�$V?8�� ͜WQ�5EU$5!d�Cdpx`sjWQ&>WጀX�O!!��?�(���+uW����t�Y��/c����K7k��9�3��8��)�m�R�R�����-Xf�����Z=EV���}�j�ԇ�@G��!����� ����h O�8�����kD'ե3��#B��1�!~���o�L���^E�XZm���������G��#C
�K�'΄�t�8��rg+�M�-蒚8#��������٬lM"[���H%\��U~���a}ǭ#�1b(�X��q��;�Gl7����z�,，/q��N~1H��d�Z�2
ш{)/:�Q0<����2ێ5 ;�7�!�!>��xAp���)Z���&��~�]����Ed.��J��K�ʍM�z1K#"Fq/w�N�Ñ�P	����!���/�{�10�Jq�[rd���xTĘ�\��c����$\ vWy�����/�(Z�;%0��"Z>�ٯde+���V����1�sSL�3)�/�>�<5��VA���a$D���CF�;K�%�fE�֑wi���n2/�1�}�ȧ4��ŀ���<�`r1g�e}9�������&��vP��@]�-s��{�Ҕb��eZ��蒄 �	Y%~KjCZ���;���;>���������r2I�4�$�m���[{�\���\�ȥ#I���i��V�P�2�|�v��y�� a.4��y#��J�"dBI!T�`n��Is=�dF�6k�\	�܅;Ĺ�I'h������C�=���R8�=V;R�$9,�o�gQ\�� �()O&,+�e9ꮡ�䢩��	
�fY3��_��`D�5<=m�#�UR�aiJ���a*%%۝�Xs����6AD1"�6=���%� 0ӭD��	K���C���8i�Z�ANHݯE�'���{�ߛ5;�Gի~��/	�׆Twf��ikd`��gX*�T���0ɟx�T3� �7�d�@�X�ay0&"mt��t���o|0<سLk2�6�p��To�ؿ Y�P&{��j�7�G�xq�[Ά�=�BNm������KgpR �0�Q̑�]s�}����W��B��+��k}s���h)����_�=�7揵�(�4���?�Ż �E|K}R��"���K��\t��6�W�qo4��c���y)�SK^�ʁ��ף^�Q����UrQ��
��h�0.rpo�5��Yr�]o��ߺ��E:zW��3�ލ���*q�sw����t�470*w�E��T5Q��"x�g�."��ҁ"IEko�~��JY8�>l�9���o:w'�E�.^3̟S��k5�Ub���5�e���e�����q�����+����W�o� Q���!s��m�x�t3B��wr�Î�ֆҞ=0m����b���i��$�'/�4:�������Wp��Y�cy�'� ��;�i�͎s�7����;�ڋ܅	D��<2bZ7�x�c��w�X@L���x֎P!jYF���x����~�Z�*������6�p�`�FF%�k;��N�PD]��u��ē�a��G"#����P):��+�@��p����˳t��oO�a7��Y��jIx��`(������zbS�P|�?B��m��O��ܑk~�!�<�]#Ip��ZV9�\m�6k��
+=SI�����:�i*	��SX�˸��Ҭ�74PcR��K4%���N,@��� "׹�|�GH6z>4�}�56f�+{��4�Jc����R��~��Ɩ�b�1���#�j26D+��b���k4�-('��V:TTefQj]����j��"#kwϘ;%>!�$sU*h��*��i�Ċ����w&t?�P:��	�Pd�5�6.h`�;��|H��7]�"ߺ�G�~�
):�v_ϱ�}�P�s��4T�����9dQ�Ng5Z�z��ʞ ʼ%,8�K��W�U��Q���&��"Oކ����N�􂛐�D#�5[hX�"\u���
s���>�}�=����Ð jX��Ws���o\�����8�4�GoN�:�}�g�h��9�/�۲d�7U�i��*������
2W�K�D�M�Pޠ������T���EXvJ͎tD�q9��j?�X�T/;Ի��%Y�5�e�d@}��&t������BRU��0�U�S�B������3�+z���h�|I��%KS7�(x	ɕu���F 9Yp�f��0V�o�1��p�@$J8K��z1����F�s�Yr�W��w��q�Oݠ���M��y��~�{ �U��Q��&MN߳�/��U>���G��.���RaF�\�s��5��]�NMk�}ˏ[�U��T��=K"<Z�[��+��v�B&�(�#���5�mHG�iZ��T �T좳eHұ0�9��.G����L�H}Rk4��J��uLB�lrZ�2�}0˚�V�8�"F,}����R<%�s�&xo��P�*��Y�Y�c�?�o�  ��J��v,��{S`$e�K�M�iA^APc&���b ����V�\{��XGa^?(1�6$# ���p��u�Y���H/�NT�!�4��9�8�@�NMկ�6]Y[�zk��.�7��K@M/��
�gI �m�>�!�.��=J�����CwN���x��3�]����B�宾k�'��	O�c�rz����$V��6�!�D�vHD�Sl�m����}%���~��칥�YH��N!�/�����s'����}��{.Q�m��c��g��i�h�Ml�?÷����i9��^�����*�CMQ�H)�x�	�i�c��p�}Dùڽ˙�?Ab�)��	|�\vPz�׷F3q�~9�m-Ϛ�<*e�(7�&�"��/�P��`!�-���[�����fl��� �V����e+�f���j[���y���'����̼y>Rl�9�-6�f{o�XQt��خ��K&�j���:��7 =�rB�:h�f��'�0�o�2�kЖ�E@�JC�K��m9Т���5{��R7�er�c�e�^�Tؾ`m%��\� [65xZ�i�2H�̶��Uگ�=.�ƶE����Ls���{%m?��~$j6�x3�!o��]���+��#o"��
O�Ш�Ϫ����r�BzY�CΖSDav-⦬�j�6���L����������i��.���C�W	��v�5$ǆ�`ا�c*=J�㿽a>a�͍���x�=bB�g��G�c�' ��l�/b+�H�������k��������wYs�(Ӧ�wXh�vV1(��RpgmQ�v����j�t��e��~&��!0�yb��=��6�,Hqg���^�N�GEn���c~'`���1�S=ڻS��L##�玫�q2Nh���:��m�Q�����+z۷��u��;)#��H�ғ)
דP�����1<$�Hv��?$Q�<`2�Y�i�Yt#��Se.����#/�a�'!�9@<�ɑ���ǡö {5��J冀����ڽ����}�s��(n�]�z9dq��ҧ��=$rKL�JY4�x~یys�]o�9;:۫�B�����;~�_�2���H0�!������)� ǱK���U����y-;�is�U�e[1���a���(�lx2��Oѽp�*;�ڽ�_~�Y��P@��΂����{����[�����������+�6}���lV7_�E�Z.��9RL���:�������)������]��kYΜ����տ9\�Z���5�n�UkX�.j��l��m�Ҫ%Oj(����_K?킞]��?���2"�U��;e�1�0lZۢ�ho~� ^��z5�F�tV�	/dS@�� �f�;:������+'�)��w/ �`C�Q.'������|�3�K�51��G�����0��s2����䛟�:�a.�sl�OgL�'	!���]+���("\�m(��xs��� ��)ʇu������>3<
�xH�SU
�<X�n�\:�t���&ʄX��¿L�ͼ��j89��\V𲽶3|�ڈ�(���=XK��������%fI�GD��,��նt��3*�b��C^\l+�r:O3��~=u��OY%L*='��>L>Fג��,>Uf��e>�<�M%U<����M��/hG~Yvi&c��E~�x��5e3���I�C������	 �ܸ�R�ͥE��G�^�����p��I&�flY�X��[£_����W0�.����"��ɛ��<�Nm�E_���"cEC�X�;� �,)e�Z�2�j�R��@\���%���O���%�zڀ�g��y@�;���3�`cvh�gIS�F�wa� H��u�����铕�b1lw�N/�������vSHrك��yp�YY1���tZ��e�B��y�R�rؖf�::S���^�ؗ��znS�2��[����N*��}��T�k+�b�R�^r�>��3g9	daiy������� i�X�5M��Xi0^�8�`��=�ٚ i�$v�'|Ƕ��|%?��s�E]U�n�$���ߔ�g�"*��*��,}� ��zc�z��'�}AE{�#���t�#��g��]�.?�pD�����3���s�IyRK����j?�$���.�FtS-�X�p�?�+�a��z�rD��=  �N�%Z�j�H҂�?�D��	��(y-�%g��%�&��M�~��7�7�Z,ދ�3�� ���q���+�K2���:��ºs��9�T�?6p&�+�#��zρ�W��n1y�"@WE�����&��0�S-$.p��P;l�-Lk�d/6�R�y?�.�K���|Zu���Ż��χ������1����.�����E��Z�2�U3~1��1���� ���גhQ(,ͤ�;�<ͫ ��΂�-cH��9}�?O�/�r����Qc	:��o��Y2��^�|��b' �X�����]g�R��W�n�e�^��y���$�U2�[��B�Tgq�"�l����,c��2=�#$Ŧڡƞ�Z�ݖwR��੐���uX�n��5:�E�}���kh�{�]����%V�` �̯�h�%�8v���p����H�W$�{I���"n��5���DǱy�k2�"�f��s<��P��ڵ�;��l�AH}����<9�+�*+[kܐ�S +	I�/7��5Gt��WE��$�[���	J}<@��.OT�VdW���M�h�l@��JB4T3��O�A��oR��[]>�D��{��$�t���xO�[�]�{x�pNB�9H����.���W))p���:�%.1-�k�4Ȍ��i�dqeLM�q���n�ີGʫc�������P���9�3�2K�<Fb��{-w&��7�@zGH65������9<9C5�MΓG���)�H���_^`&H��w��Á�u#�����@��>N����j�V�X�l��?���:u5f bM�6�5S ���v\���Ω$7��]6� ����˱S���;��Y�b��SE|���mY�ؼN�|q�PC�ui�o^!6C1t��r܋�6�d��*~���)i]����%6{��Y�p�	lw����0=;�2G���(b�z��{���n~�rBn�G�?�.�Pp������W8 �*���ٷ�\����~,�%�7�8ڨ�L�{[l�d�{ԖqHd���&���}�}�ZN'v��j��"J�eE���G�Br�W�Xt���>�rP�/$����D���"K�#�z��"f3PM�㛜~�Y�^SJ�74��#�h�0S�R^ڜ�Uj���]TI�,�vhJ�?������r<T<Q]�5d1
�p��]�dN�?!���^�{վ��V�.(6x&��V<Aȉ]'�j��f���W��3�$fB]��o*�Ѥ�g���&�,�'^~���껹�ڝ(��s O({���";c1��}�=
\"&u��Ѧ=�`Z'�����L�Ą �^�@3��r���S��Ѓ-�Wc-�]>��.4T���Ja��r�TL(�N�q�P��S�:k~>W�Џ/V��k�<q#��ONd�t+������vZ�2�Q�2��""+�OӬU$|���O�nbE�1���o�T�j��̷;����f��g��=Ū�Qm:W��;jߓ�3���)WJ�5Ί�0y��%�Mo ;E�b�CW1]x{��a�N�Dy��;{=�ֿJq>r>:�Ņ��2���j/9�����Ac�����9�Ȳ����+A}�k��a2������L%���h�ᾳ;1*ў�c��n�Qϗ�n_b���-��*w���z�|U%��ASE�Z�ro�/�1�~��f:��,!�K>{�gTT!�&��E!�A#ׄ]���K�ҜH}�l<O��q��K[��T��H� 07����'�/����Q~�4�=�Ȉ#���ŷ�z��Wt6�P��V/�U䲽z5|5a��Y]\D����ia�	`�IxQqs��#E#�A��QrK�<�����"{l�\��\t���J�ۗ
�ѧ� �zB��y��ǂ�/����?G$KI7���b�e*����KD�>�g�5�,�����G3��ihS�T��Cjt덒Q��m6+��|t�o"_I�K�H%�g��+l�ӄ���t�k�?^*���3=4�[���,�0�9�mx9�؆
�C|w�8�޳O#sW��Q)���[�*i�o���aZ:�ۍ���ʚ���M`�z���F���cb�� ��P�y,��� {�:�!��轖E�SF�89���ў&=_�͚��x��|��	S�Y�0
���[�� ��=��.����x��:�i������DI�36��/���9v�@�$�8�כ�:߷͓�?V�*�q6��9@�Y�ȇ�0u��2����/L�o��=��Z=��;�+A���+����8I6��>/�g�^HT^����������M��l�'C%e M�y�Q��]�� �+PQ3y���F8�m�� ��a��G�)&D�u�W�+
x��z]�2Ɉs�s�XI5���/�aؐEB�(���c0��r�;��6�&�E�t��o�T�8B������M.�8y����z:��z~�#�O\���$�s�{q�qN� |��]�IL�O ��bSc�u���o���[���zI<��TjC`�]�-6�w��}b���	+1���¼��[�w��)����W��O�Pi�5e�u��uq��#[T/wd�^�w�4�7j �?��5����r�4|���߬�t�M��3�W2�pu�~�8���HI����1���^͗\d^ ��#���~�� 6����И�$��g�tO��v��d���U���6�*8v������g�g�:��/=jL��/+@,l>k���V���Ĝ�,~�`����h���iy&䆎��n��=���A��	XE�_�ϼ4M�zL�|���Q	G�6�{��Wg�r�b}�~=���yb�/E�]���%3f4ֳ��Fˎ{��0)n�o�V��f���@
.7y����5U�Z������咲��."��ʈ�������b|����+,i%���<�-�wb��c\l��jM��`_Z�`-k�1��C�D���{������;	t��s2^�2�n�f�:f��!��(�8�� �{��"�p�w�7lQ�h�TŒ���q����e�n�C�yY�\y�
��mn��!鴄;�l�2]�A������~��躖{�RO2p�j���H�|h_/�>V���܉.�}�B���z'Ai�'����P�ȑ�$��o���O_��7����$�T�McU�Q�/|�-/�v��5}YS3�[[ڶ$�Bn���>�I�BP��@\�A|�OU�s}�V�w�LxL%�>�_��K�]��Q���v�CQ�G�UK�Fv����U�g	�ğ��8��G����� Cd�nsN%'H�q�h�Y���G�ĥj>u�1��Q�oCY����ך�!�L������c��$�.��0�4�8w���jS K֝,TɊBLW1���0�Y���<���[�>}<\�J�yB%Z���`�$R���C�}�yj������X�.Xj#���{z�v��6�e99K&b;��/�!~lR�|��@{-�}�Ƥ8f�5�f��]u5��0VB�V�;%�f�%�� S�q����Q���-�tˤ���8� �z)-n�z�ڠ���X:���7dL�x*"o�ov�9=���Z�d,-_=��C�J��R�;4���fϱ����\w_a��L��}.�F(9�,��y ���k�lW&��}|�hVΤ�*Ii"
�JM:��_�m�q���_�������h����&�D"	���5[:�ը�'l�Ũ|�\:'c+(@2�fE����eB>�-@CFI$|N�sn�D��!��Q�	��w���"��ډ?��+��>����n��#�"GW3��m�; �vuL���P� ��T�b�6	�`�=����.Cc<�>��ޢ3�'��k�q�l���`�]�%,���mL��͊�D��dl)FY����P �a[Y#�^��9�]PE������JD}��	Fγ�M����g��ϰ�vB��?�Ϋt�Wv2����bI?�B�b<�\'�|I|��T�"������iyA�� �0�y��!V�"V�O���8sǪ�l�:�ܥ�,*�������u���5N�����f=9a� �i��$�o7gg�M�MѺg��+�)aL���K�R럠PQقa���	;�V�w�Zˑ��<"�|��"�k��I�./w��S�`�����إ���M��`Mȿ�������j��H�v1#ORw�D�0Ԅ����HpLs3~6q��O���<��=� ٪�����g$�vʘ$��G��9��x��vM�5V���>�G��M<�:�f�+Y `�dV��!�^)$8	88D}`����	�s���X�t��
�<rayԶ�g������דL�U��ݦ�ޡ*��F����v7�I�P�5��R�<6��m?��s�ݒY���ꋬs@��]���q��	��y���>o����
f�[��+��������h�D|՟�l������7k&#�G��>�Mz��T���A,�:�����zpjP����Z�j�6�FT���4�� ��,�q��ϳ�{G�:�J|.v���滘u�D�ϤH��&Q����[m��#.��q5�Y�5F@!*^S��ܬM?3�N�Q�#��?Z�`!PA�y{����$q�y4d+��X����k6�>�=�Ͽ<���6�9J���<�tM,�kՌ�nEw����K�q6��|�xÐr�S�mB��t�lӼvX�i���E�4��dAQr7��{GBI���������L�J�.P��{s�xT��z���o���%����o��i� �-#H��h8�)�/�����EgQEB)p{Ge���'O��um��@^W����=��╃���Қ��a�\Ӊ(:�煂uJF��^�3l�n���$ P\W��/����L��chmPs��<�P�#��D�F�\��m�YI)�@bda��.zw��g�	�z ��"�\���Jy6٫j�A�F� �ң�p��F_�gj�{kQ<�P&z*�]�}/����t�����"LҼv"��V1״��L`>�s]{ -/r}�MUD��;��묜z�A��O?9��Bӆ@ �A�'�:<
�P9"x���Q%O��Ɣaϯ;򜝊�RZ@�h��e�޺2�C���~�(��r)�?���]���m����C$sE���N�	\x]m��ѻ�$�C���i�����/7/>�f$	�p������寃ИC?!�o#���V�=j�CDZh�� �4lM��e��?��M�o!X�W�� �Đ���"�8�X���M?ъ���Q�BQ����'Y��L��O ��[il�1,`��������������d}ٴ��W �2x�Ocj�5iYSs�߄���f����D;Ɗ�Hn%�:���/� �I�q�K�Ñ��Ox�݌���n����6��5��|���_�
��<������\��p��%��~n��Vq0�E�T��j��1��6�r�X��g�G]VJ�U���<��7�M���}u3L�sU}#?K˧�-"5�,M�x�3��\Yܜ:��j���%��l���K��r�G���6E8P'w$ԟ��k�.�TONL�e�v�.^�mߢ��0x�K����f9=y&�7W��� 1�{��r���N��J�T&�A�g�Ė��*��,}�L�
��'/�?|�t؀n
M�؋g��y����2�ۡ]�ċݚ�Zj6ǩD��������\���"��#!a^}�Ѩڹ��E	:ѾW�X:�;��-â��{o�x�#��`��K�6I��3�Q�eo�v����2�CRL|C��c���K�����P�'ŕ4m���C ���*�@>h��Zj�`~�
���U�!t�G�+���9v�릴�¡����J�;�����q�s4)����	vzY��ZP��+��d�2������G|N�������0.D�?�*���hgbP�y�ЮvX��[[�2�׻hX�b��c��᧤��2��  iLr�h�"�;���K�LśPF/���5@�:֭Aq�?�U��Z��f��%��g↕*C20���=ي�=6(<5&�y�r���%4A������	{;2o'���C۾�R��-��gM��Zy��7O���BVRG-u��Yy���P�L�j��-�C��u�l(`aa1|(!~[�჋�JrGm����#S-���:�v
w����(Ld"�������zz���G[ln%�nWgB��qYJ�V�؎@G��%c{o^�Z�8Wꓬw�R01ӗ���N���o�qAF��+YO�<�oo�HRJ38�GP�Q�4��~_cU�A���*��GE�	t��̾|vY��:��0=�q�2��d�v�Eٵ�t3-��j�P�:ry�L�`B��Ѓ9M_�,G> �\�4�,7�Be���$�a+�"��胮mG7XI�Lp��0��iE�-�i�\����F�Qx�o��K~��So�V�/������6�C{-�~�F�7wF(���3���Ocm	G�Q!~aL���} �|
~Fzü��ꌵD���vn�0�(tAW��UP�T��'�mwz`�!:����	\�9�üjWX�r�O�n�6C����_��^ci���b���M���j�U�Ao}��������z"��ps$i��*ia��.7.�S��M�	�s��$����&^Ax��n��������;�P�]%/�LWy�fF��{cF�epf�����t�^8)/�b����#�c���&TƋ�Ŭ��Ӥ��>�K'�1xdޯ<8W�?� ݚ��Y�Yg"�#��v�Q��_��������ޏVk(_J��^D�(�%���c��������O���5s���n1��/��F췪��&i ��h?��$�*A��bQ���e9�+�f�%�A~2)�4��$��S�.W��~��B��*YM��B쵙���I��ܲ�6�Lze��5[R��U�<��^��w�g���=q���h&5>�}h��s�x{���+u�t
�c���*E(��&y�Td� �=��U�Ƴ)����Ը�R���d�u�Q�f��߂��T_�q�U��G�
f@�>b��#�i�wM�F�g��\�#��^NU��o�6;�b��^f$���ȩzOc��+j��K�B�)}�\����k:=��ey'��t��`#�	�;	B$�b�r�D9w�b�*�/�Ņ`����˓`vĊZ�q(w�ϥ��X�`:S�����a�b��SC�Q�.��X!���T:c��t�M�T�K��I.OZd�WLR˄����c��D���U�(����T�$�oJ+����D��MX�kM���~hM�Ն�6!f��9�*wu3v����G�Rkb$�P�L�f�����m���X�E�mA�.y�ޣp��
�]�j@(���1����{��g2;��D��q��6�u O�i�0}b�&�['ҙ�jd��9']Z!�4Dl��4�����d7�Z}W�����n���br��4��8�P��	N;��v�nu�{y�$9�uu[gf7O���*�c�C�aG�B���5��YǾ6���[��e�ˤ�8:��>"0O�I���G���u��W-��+u��/�n��[
���O��;?�wQ,V[�ڢ�֦��݌�!���GI	�A����(��ʪԟl,�-���=^&07r.w~���
Ж�;s8ea.��(�MUQ%I���Uv��7���9��* �&f�P��Ĥj�RoF�ք�l��Z�m: ����Sa�")@����������Y���C)%ԴF�. �O�{��ɪq�����D/�(!������/.�@b)�`#�PU|iJ�d�*���h��E��nI�u6�R���/8k����jl�/��9�*���)=��=X�͠� ���MXMM;8>[�|���z��f��7���4��{� �B���OeUv��@r�_�������kV����^ІNz�d54z�Y�.mQ��}��F][Z�Z[be<����e��.z�������?�����R�'P�aǂ\8�+T����B�]�h��|���!����m��.����/��f�qǎhF�\���3X?1���h~B�%��X���b�e-<?>�� � ������'4a���A���+Zk�&;4p�t�Bl�}	Y��٨1���RB@Iن�K�
�e�f(���H p=�LG��]����V }IA2/��L#
D����J�[�D+�@��v�׎+%>�ď�q��	\cpn6����og�<KC�?�e�D����5�΅NA���'�^��os���8�߽E�ђ���Ym�|͂��z[6�����+��>�鏜u8�D�X�uq-e]�L�-��.��а��jl������L�j�m�=(��ë��̐��-�#ɽ��vs�5�@뭠�m��|�_N�88h�	,���sѲ�A�1�VdT��ȶ�G"���^�Ԛ��ě��W�2Ͻ�#�ˏ�z��b��0�jHt|pVu�E��%o+���k�Y��ܿ��k�k�o�`��T��7���H���s�Cl�{n�+��ā\�O��Ě�2\ϐ����f�T � X�Q��?�&���f���`�#�_�ˆ+�c�2�4��h|\J
��z>�@q۞l�NAs��2ȋZ
��y��)�䟮�u��T����tNFjwv�
,���»��M]���B{��?I����=�CNت����J���x+t�x�_K�Z�!h�.a����۲�I�
��r�oj�"*n��R��k=���3$��sL׾>��d�$�pwK�����,��B3���o���3��@�l�&O����O��g��$� ��᷀��d	4�A���|T���0<q
�r�h��a�����e嘯�d���^��_��:Q�U�Jש!�چ�T*�N8��5�`!�gM�%M:�ڨ��4�ß�l�f�>�m����,��`��
nf�e��߭���Q���s8�(T��pt;�Q� e���j?����-�8G��:&�ݹ�v���6et6������w&d��x��cl���'A<�X��l`IW-A8�@��1k����\Y�0G�rl�
�ꊗ'�ȃ�(fO�DON��<6@$�fo�W�Ʊ��A]�&le���i��v��nS��F�K�<��pH��rEh(���D`����B|�''��ӵFk֒���_¿�w��Dh֧�Z��s}�+�Gڳ$krn����j@,�;�y���1[�������$� "o�X�*�Ù�t ����h���I<�P�^Q�ܝ��1&]s�W��E�h�n�fkع���>��x'���8��1����4k���&��o:\V����A�	�uȪ�������j���L�칯e��b�c���{�G8��r��)��ڕ��:��}��>&Ҍ�|�����C�&')혇�j-��rȭ'�:A���k���^��bmq%�ӚL�`��]�X�S��`�Y�3R}�v!?&�T]�xGg�^�U�"6Ļe�^��^����,��g��Hv\M�S�_��Ge��3:�ƛ߆#�1#9D���)��E���E�K�+��ؑ3w�|br���a��Dћ#�ȁ�B|�fR9ݱ �TU � ��f��H.�h�}�Ƅ��r+�yM�݄Ă>z�gj�i��"��:%i�3Ɩ>��H��F��~_�Q�J����� y�$�7���h\$Q@�l�,��
/W��<C��Â/2�%׋.��G	U�*�f4t!�)Cxf7xĤw[��lB��3�mY�xHe�k/�ÿ׊YCG8�0�
��D)�������4$��-⿨<���c�(��~�QT�@����Y��?J�y	'�o�P��Ig�S��N����K�X/���(��VMﻨ��.���]��6>���;t����L���u�1�ݵT�w@�Kژ|Z�"x1/��f�E��� �:�%S�W��%�q8�����<��Ǟ�A�w	��!çb9�ؗ��W��ѿ	�+Fs�q���O��l�Pl�c���p�f�`���.Mʢ����T�j)*~�4�F�i��vC�ȑ&+���-�hF��hS�GG!:y�e�d���\�2��	�� ��͠����m��K�Mm�Z7����$�⍨�8��GQ�b[��t�r�4��3��$zWP�}SGm���Җ.<�j �����H��J�裾��%�>�T������O��	��i`A~�k���`.�Vި���?MA`|b��^����݆�w������;���;�H��)�^%h?d���l�P�tL(��]����	�k�b`ߙ��_]�ړŋ�?�(���6��r��#2٘���E�b�Nkg��b�����r��b@�D�z���׌�9��3m�˥�_	R|	os�x�y�)v*��Jȃ����*�V�Q��e��:#�2�o�Z}XLiY*z���s�gs_�JJ��tx�O_�t'�i�%�lZe`Z��&5��$�&ߤ�%{t
����ɛ'�#M�Q�sB*nI|j!��:�	!u��q�^���}�x�2�݃Y����A!k%�EO����ro�J�ʹ��XB�`�v�t(��!�Hx��sTYH\')
o9J�����*�4�ʄ�Ty��U�Ζ��t�v��|b�P���Ja	���`w����P�O�u��m�LX�}z*
��s����o���1"r�?�E��������P��QQ%����3�Kԭ�hR�����E8}|f��ի������?��~��#�^��VI�-6�|FĚ�~m{PH����c+\�S������:Du`��L�GJ'65�z�/�\q1��{�+y�U�2�ñ7�w�\ڬ2�_-�*P�A	�KԬ�ٿp���
��`�4��MX5�ND�����ѱ�Rwv�:�&;lx��=�(���:���.�	T8���HS�q��mLƛ�'"H��?�w��.jU��*O��@��E����й�d���
o�s���bF�Og�I$FbK�0]�Y�c��g�?I��g��
�����
=(Y�U��^.�����������`pQa��j��e1�?��mz/��� Ī������y$[�|HY���{z�VR�G�C	"�����ō0#�Bq�a��퍪n��K^�q� e�C��[�q,�K����0t�V��HQ��ՙb��x�{�u�-��ga�����T�J'a{K�nK+�i�i��o �=(u���\|b�ޡ��W�%l��<(ɬdי\1���L~�6�4a�%w�n��o�{�n�"�b̟��Y��]�n~���@��n������7����8�����~�<A�%x�D9W�2I�#,��-I�n�Ws��M���-L�iq�ۏ؝��F��.�lec�c 2T{�l<�t�!!�>{r[�j���1Q��4��ǻ{Wq|!���������,G�J-��E�P���l�Wt�]r0��+(w8ʣ�[;��oRHq��� '�*#%W�D�f-��C����|�����x17�k
P���`�?����p���_�;�{�:{W[MkNQ��Z[+���_�bS c��v����"�論�p����HF>�]������uvSnrq��`	�m�c@��NfKG24������_r2`��V�b�'>�E0��ǹDu�
L��:�q`��=x͆'�v�"��!V�~� (�v7O����^`c]�"��S�f��ZBs�L�7�gVf��r�S��c�֓ؓk�U�l	�12%���6Rq2���T9gR'��R���%L��8�H����(�<�.;����%WG�㺏{��t����S*��t���o^1�m;X/��U��$*���̑�l_IR����r����ǜ�=m
�W���f�S?񓤛dX:����+%���I��~/�>p-��.��zΟ�g���-�$�#<�bزa�K(�B8^�6*F*�Y��I#�S�uA�[�����X����׫���Vb^Yly��̀�v��~p�D�EI:nz��@āQb�x5�?@�,���gO��N4>����x��rO2��ã��h���j�5�瞋\���iK`��(ã(�F�;�T�:�b�;/os��`h�bz�MI��kCQ�5��zp�6�� 8�pθ������Ϙ-ܝ���kPa!Y�S�x�FV+�GA�m��G�	)�#�vQv�0#&(�sN�s(�%�G�Ġ���q�*��g��=ųd&˙3{�FX�Ҍ�'I���R>9�u��;�а��r�_���ҕV�f��A�����H�)��]�,�k�9jm�!��M�9���,kO��?�u�D�ֵ�$�q$��W��������� ��K���8���u6���[�����9<\\F`Ad�(�j�N�P}�+�-&5���x�e/�7�ǒ�9��(���x;*�o�t�U�
FV69"Wp�&��'A��(E�qLՅ�����s&���ꅄ�	ӆuP ��m���}I8֦5�/'���M�NF�/+�(:�)� yBȹ��v��G��o�8YR�XG�V��	�d����e!�	��v��p�yc�xA��@] RZr�	��	���	܋�̋p*����]��cKZ�2k{��8;R�0u}4Q�����V'�?~u�L�lw�y�� �S(�?1����é7�b<~�}�ƅ�_�qՑ�UA��\Y�R�]ɘ�ڮ_�L�&��gc8�W�)��(��Ldj��1f��93�e?�&�7]j#� m������B7<I�3�U�6J_�C7�^�6#��xO]S��w*����̡�6� �� �K�(�`��B�M �	�p����SGT4�v2��	�H������k��NOm,&��8��5Z.�����x�I�=�#yQ���}i������g`���c[C�D]�W��	ܭ�-W�b�b*�i����	�^)�uп�!]�X/r�� ��
��\�+��ِU|�9I��c��<�P�f���Y;����A��g�i����6����B,��@�-�&KZ{Y�����2�����E�]A�?�W�&k<�.*����Eq[,v|�db����������`��:�jK5=)��7	�"��W���loD�N�+H��c� avrb��͙�[��̪ m�^kM>����P�HùpZ�����;ґ{ тv�&���Fvz>άJ?O`C
�#��������~gP|���(��5}�F�|�<b�;�wAʝUQ*�8�.�|�7	�(&��B�!���_ӕ?S�ru��{?���2F�I����k
�I�*�D�B�M&9:�=&g��c��'���k��P[�\M����8@;ߜ�[��ƙ�Y�t-PɄ��X�0�CX���:^������y���'v�x�0!Ie%�^z�)��������T|�㜳 �[��j/���H��x��B4v���4?�Y�,x�m	[UlѨ���t}3�TG1ϗ޻P )P���B�#!��p�,��kkp=�W���]>�����!�a��i��#�_�9^�qb�"�d4�/�-� �(��<������<�E2+BrK��E�ﮊ,�ۼ9޴�|p��pj�*�m��Vv�E���Z��6��}��ɐ&y~�K�N�@�@ihe��X�e/��y�$r=V�+P�@��$/��&�}U��Kd�Ϛv��Q�4�.�/�a�`8$����d�{�&&�;<RBU���АH�c�<>!DM��d:{���iq�=��>���E�	j�sd�HPԍ*���f0Y��3��l��Q�Zny�'�=0���}(dS�w�><��`Q�#���HDLv��3���d�ш��&m��{���۔���#�y/�e�HEU����Aڍ�2n>�'�H�#�:�t!�Ȅ�bt���a�`�IC^�5;��K�!���h��Y�LDd��`�]�J ZiO�*�I��@j���r��6�t*���q"=W�T]���r�W��8Պ�m%�g��'Y�Tz��(��.z$�t$G$S�|�?Yf���#�q�S��@�G$-<������Ŀg�U��<g!T�4D�J�R�i����\3!:6)΋Dd��g^9i����c+����?�E��=iD�`�-8�䐍_�3��>�t*U�l6>��з�O���~�L�#�k��V<�;�ZH�
;�]G햃�>�f�� _�{�4Q��j�*o���(?�?=���j��YJ�ԡ��z׶@�\r�9�t��-�}|�;�%6�����@T9Oa!�8,��л�=}�8�ei%���wƁ�r&�qʽ���1��xE�p� �ub��(����&p`�@�쉬�@ᇅZV%�6��s���^�W�o���v�h�U���t��3�2x�sD�Y�n�Z����t+|��ٰ'g��̙
s�<Z����]��+�w^0������8Y(ܹoQ����ɖ�X��Kr�G��(|<�Df��&�������_~�l#8��>qqc���>_���cy� ����ƈb�ࠧ��Z�:����f�Rt��,�zȄ�K?�F�K��_��d^$�"�����*e9���$��(��\ZX�̷2s���_H����L��;�L�Hw����8���/n^����GEP]�guwX`�@8/�Ґ��{Q8T��+���j�����n��tUMd�Q�my/b�:��,�Sd)ޫY���8Ow�{��ˊ�'�X���w\!�Y�s�e����/��n�&G��K�i��E����lD���^�B^����w���b3�Q��� ��ٗ��@����;6Ֆ��T��$�c��tx�U�w��i�+iE�=�F�F�tXO5�\��W��#�yYͪO�t"~�o�F�rU��
�^��܇_ӟ4�`H=����w��~s��'^mna+� ՈSq >�zm�:7P}����� �"�D���px�2��MPݬ�C�(Z@.0#p�ӭL3��i �����
u��R���9bCBk'�_l\z�[�Y ˏ�H{�����O�<s�⋽�^
y1�}AH0$�Q]��l�(�͘� ��@5A�i��H�1�>���K��U���h�����c��Z�-���帻�,��?m�c�Rl���2^�������p�����?��ɵ��.~tz �e����]��GJ���4��� �����@�8��äX��h-�t�Xhlx�����rS>��i��]�#ۤ�t�w.��*���1'�A�d���X�q��Јm�y�k�kX��İ� &���0���2���v��7z��e�H,�kB�mY��t���򰶢v���;�(�]f�la_jU����H�����:\����svUT���X��W�C�� `zԱQ��2̧�a�ᐰ���i0	�PQ�XŇVS�_c��S���F�a�ѫ�7�N�hb0�r�m�9��Ul�)a57�O1����Si��ļ;uë���e�R��yqL��Fތ�	�2ǜgQ�w�t@𑀜�g��l��o3a�|�9jr�����@6T����e��&*iCW�x�\�@��r��[)�]�WY?�_��9i.��2%�n���eb�jBMj0אnr\}_��q�����t�?�W�|�JQ��0K��5!v;�g�-�
T�\���mjp�95P����
��,Fv22LИF�0b��A̎����I5�&Po�a2
/5q��9��x}!�׬*�W~E�r���f��&���e�Iζ4�mu����]�>þ[�!��0�岞�*���Y�0`0R.5W� )-�$�/Q����9.k�0t�J��r���ݔ�,��q��z�D��z ��+L�eS�缾�����?���k=rt{��|�05\��3�a�	����TN���ox5�L�]��"g=��S��kq����^4�
���*�$:��I:DN��B?Wovb�i5�^G
{�^�Ӽ�At�r �ʘ���RDon�zP�>H��,[�S�5�e�������;� z�k�e����!�A�S�0��ZcXE}�[�x��XWTǓ���d��$�R�TP�m�,�эh�:�Q�N	���*�%/kRB��l�1�m��a�����C�w:�/����jn�M�r�E�8zΕoC��\~<��z��B�1f��q^0���łn�D��0Zgs��	�y�IQ�f�m���V����Ǚ��r[O+5��S�wU�y��+li��.�n��~�g6�e���Z����(����!Z�LrǛ�
a��16O�*^�����9
��X��V*��q�3K �[C^��1��_K\�Dk]�Ł�F��X�o�R#��R
��qsU*���ƲWy�J���s�G�*:Ǒ�1%�ף����5x?Zn�٢�U Q�P-`%jD�.Ї9��B��آ��B���`M�Z�9�h�&f��i�S�7Y��7�2=Dϭe��N?�1�"	_�/�h�^-1h����f�>3�	�Cg�s���`m�s�W�pෂ���Sl&��c�ކ38SV �Mk�6��$�o�#�r�YV�z>����s�.H���]���v��e��}5�HbD9
�Y{K��X|��z�n�/�Z�Z�;_��%v�YpG�T��pv�5b��>��u]�d�6����mND�����@iL��J&^`�j\����7�����%�4����&���PV��|�� ?lTl���j
YKL�r�0ҿm`ˮ��"��$�T�?���;�#R���Ƅ��4tZu(Rsc
<���l��Ru"���`���f.*�ˁ�'�8�/�`��/0Z�<'y��鏅}�
f������lƘ�*���?��P���JW�*Nl��'�RU�&��&��?u��7$�4������򑜄Y:��a��z�)�+�pra�|�_\�L��q�*�H, MIG�3�2v��cVI#�'�ʵ��c��jtG{���`&yi�oΰ<2�ei^ML��c}贜3�
 '�$hE�%T
�4ҵ�a �K��F��!��5���T7W�gF,d�9�\�u��:*���c�p63�T�UVS}�ޏ����I590C�*��u�Ո�<� �g�
(��¦���nڻL�tU����%�^��Ҙ�낟�W0�|��x�ʮ�En���$�#jǨ*��r,���ƌz��,�" ʙŅ|�ǸG{�s��R(�_��A��L���yC�u>w#��t�ú��r���v�1j�k��c�cz/��ׯ��B��Ԁ��j�<��Q�
��d��_���������	��Ɣ��.��^�mF�	͟q!]��I~��'}-��w����b�o���oh��xX9�/�F,��ׄa����9�4��SL{�

4?k־!��*������j���Cv�������;؄����f!z�KE���.��#\��X����8P�C�@�7�������<���.���)$�o^��]�P4˦��9[��iz����qc�'|d��;�%9��Guxg�RH( ��e����VH��[K��ЁOe�a�ÿ��<� �?��/,�,q�:Q�mN<���8%�T��N�A/�*��X�b�@5<�oh���_��o�&�Ez�1�y����;?����`��[�%�P�A���K�7Z�Q�sX0�퐶����q���W9��fbkg��0q�X�'���\��-����yZZ>����xȅ\<q�f!cXT򌗓�*�`%hQU�r��{=Xt�C���q�ڦc=TKz_�-�y\������F�Dq8�Z+�1*���m������7/����F�Y08}s^[��Z�$EU�)��vPl����%� ���"�Ȝ�7��qǧw5�� '��zL�>�������so�4�A��,� �miH�a%�%ɕht��\j.Z����R��T�Ӿi�,� }B������;ژ�P�5qnf�*Z�w�b����Pq�#�ԩx�Q{m>�qǀ�n���mT�( ��a��T�>�٦ /�m����y�I�
E��RW7ǜ�������`))�\��H�zc���b��Bt,)M����-�4;��)u.t�{��W��=Kb,Yeh�����)��57�a�F׫Sd�x��Q,���t��9��D����D	w-�'�,x�ǌj�-�����s[�U=�;�~d�ՠt��ǻk�w�h�=�xM�.��Z����/Eas�'��f�w��m���3oؼ��7:�#�s�����LM�n� )*.h�[�+�>Qx@��~�����6�����xT�6���t��i  Jb!ֺ��]cֶ|��x�^�q~��iC�c�}+�.�:�M������)�mnnؘ���b����e	�2e��Y�rv<IZ����s��y>�d:cL�W(h�rG�n&ĕ_�%6ƌ��NS�g�^��6��)�%D��`jx�$]JY�c�lǗ�x�<1L�f�֏L�bf�g���o��MvNl$X<�O[����t���"F#}��fk�f������i,6��%N�����+�`���q$���h�q�8[2]�����*�p�V�l��]G�ӽ���}�wP60̰�VU�K��q��������XXA�~苖��,�f0aGAE����خJj�V:Ш���g�Z��:n=�T��6ռ�M{��5��>�����5��X�"������lR�[Zd�!ڌ��\����W)&\�4�F�p�ojh�l����H���^�@5����e���Z�x��|�h1�n|Fs/�[��h�Y����o+�ݢ��<��I�0[ݠ.���;j�C"��/m�e�x��ؓk-'��tp���*s�bʠޏa%��vA���h۶�Sw	�B��-�_jՍ�C7C��\�Gi�&ؾ�'��`]�,�z�WL[1Y PQѐM޶�M�X�q�x�	�K���꬯���^F�X4R�*")�l�y
3���n$��F�Zl�șb ��;�)����J��OU&���kܼʴ�{�0�1z0��/���$��x�V�*�;��5K� >(ԟ؇��5��Ϭ��V��a���e2�<v8.V��7�9�J'0��4R���`�Ev���0��G��өј��`E.~��i3_'���cv;�;(���[&�e��c�df}=��a�����	�6i��w��i�ѓ3._���()��
]C�o,��$ɥ?��ު;v����k��2_�k14��Y�@�91��4�Z���+T�7$���FfhͿ-5�Ȥ_���s�C�"��'=Vw!�b>B���$\}%=��gBC>�·I�P�ы}�-��� �9\g�/@�m����U*KD�T�- ��P������Wg�����Q�4_�0�fe���ͤ�r�����h�����r52��ý��q��-����9��640���`�W�h�i���a?c�ej倨��]�9N$lsY͕���ǌ,����˙��7�zgә50��ӛ?\s���XݶF���Qi[ez�C�rL�����}j־�r��>��匦6����7n�{� L�گ/ZN�啹��o�b�椠��6�W໕�	k�v#ĸem��ɮ���9�W�v�g��!?k��
�D���7c����
��⛒�#��g�n����A�_�Ȝ~�+���Ӹ
��9đ(��^3��|�O�~H��,g�&g�_B��B1��n���x�O+��8��<�jw��G���������l޾_�u]]08�	��v�!����!��_�� ��:��#��*m�D>0/�b�+���b�P�O'wY��I�>ނ+���[r���J�f��jRv������8�Dh�_�I^����9�ht�_�����яm����~��M�y��6�,��̦��o�տ�gaT;l��oe\�&K��k~4�	P&Bսބ��!.��D���Hē���XA����9?��j��9���c	��<h��3�I>��
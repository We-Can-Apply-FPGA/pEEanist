��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i��������쀞L̓"�oܜf�~�5@�g4�5�	�
����,aeH>)�3+,���KԾ�D�X��x���ark��!��H�ҫC��\���!Q{���,�1��؜�C^�D�{b�؏HltH�F�X%dAm\��k��4H���5��p@���9:0�pȫ�IJQw�	@l}NT�{���r)�w����D(1( �ް#ZK|-V��$j#�C�h��U�*��`�������$+}�1Mp�V��K#�� ���rȗ�|�X�9���.cX�s^�_��P(�p��y�%�`��S�
�o
����lhV�qe����
�8V�K>.�w`��O�C�1f��� 4���T�Jm�(Y�z��u^��H6����~')�Fxe��
�f�Qz�������8�3�[��E]�A.�F���J�x`O�KV;d���3�|�B~�>Uh&�!d�v	u�o�����C��ǈ�x����Ѣr5>Y�,Y/�$q�>�(��}�̞�m$�]�������H�Gs�pVEׇ#%֮��d	b�{�d~�d�v�3�X��=O���d�\;�͢����g��cd�c>8�&��K��a�/4v�E���N�����bͻ8~cx$<8a
�VP�߻�6�o�b������)A,������1ğ��yE03M~sU�Fa&w��<�� ��V-}X��S[2��͛ޭu�E"�����<�3����*����K��½��ع����}�rd�s��!h��X����@c�ݖ ��`��F�x?�#m�L���C��P	]���"sK<bt&)@{`�@>��B�0�3������&��L�o�d�f��p�'&��i`I�����Ʈ{��j�9T�����o�	��4��+��gh�e��6�0xZC{�m4���_�.1��N ~�� �It����<�kMF٪�I��3@?��W�����O�nVnM ������Iˌ��0@нn�g�4-{��/��s�ؕ�=�T�oJ��,��Hn<�,mw�#����Q��_҄|�	���x�x����g�@���%�S{)V�4�w:�)��jjF0}"LLU�j�21�,�fy=��V=4�;���O��|~ Ui]�X���m^sN����y� ��˧;�: s�?�0��5�#��GŞS���+�*���M"��Z��!o���F;.e���!aqF�����M-���o�o��Ĕ��m�P�Y�Y��f�X΍h�����ղIIfX�G�{�k�0�`����=�r.����F"Q/o!8��%vc�09N������N����ErU��	r�cD�:�N��q�D�ɩ����)g�o�?�4�EjNg����dea�Z�o�Ġ�m��T���Jf�0�Hu�>O2P�W��lS ��>:fIw�By��x�Ŭi_!`���|�1ַ�v��bo�$����)f�C1�N4�,aI]��\��B��p��L�}��(Em��?�ś�̒�l�NqZB�ޔ����i�A@ƹy����U̕z͈�� �A^�'��Re1*�W�����#5�?_KioKkoѬ@O2u�N�{��P����Y��#��p�S0^�ජ�Y�	��h�
�c1ۼ��=�����b*-K���GչP��>/�1K�������n�u,��~3N��j|�5�B��� yCJ���|�tVףw�dI��o���Z�YKa6�B6K�p^t$���a�9�@G'�Xti�T=��Lc=.]���@åx���	W�t ��JU�2��ߕ��?�� 9@��DI�)����()u6-gy���͒����LM�0KX*A%�ӗp�v���qw�3d�$D=-l9,�OvUB�}�Zc���<D5kn�9���U>��s#5�b[�R�U'h>�&F��o�^���L��X��׸|�W��jR=��2��is�T���q�Ly��m'3��1�B�oA@_�|~�X��,�tC ��+ ���l���eaq��I�/ɵ�#}Ec�\��(E?�	Z�{@+	�-�)������k��x�7d���dD{oS�Ԩ�N!1R�^�~ D�����	.�s���;|�h�ݗ�9է��҂K.�C���u0����Qs)���h�ܮ�(I���25������Իh�������JFAN�-o=��g��O�)�	��Rh���Lz����wxa�xG%2 ��U����4n�tO�����F�;�Ĉ�<�c�'�N��B> ��1rb�Hc��W��v	q�06��?��t!��d:t{;\��$�r5�	Z���?u�;,8�9L��q�x�XG)᪝>қB5O��3���k.p]��!ω��͇����$�v�$���=]ȷY�4m���W%�=��C��c�� ���6$�����2�x�����Z�+K�N�ؚ)��}��x�L[���O� Yu^�d=����u��5�/�)����f���3���l��sW]6�sZ$�-�ݽ��3�!�7Z�0���x�G�;Ϣ"" �Ԋ"�0������ż�#�����:�+M<�}�^������SU"~	����Dբ?�*&!=ؾH^A�ʵzSG�3�������)��5�#yQ�c�ٸ\F�N	�t�Ā�Ng"ǚ��e��7p�x��D��g^���rf�z0��FӣW1Zk|�� 9����������e���쯚����@���]8���y~e�0C�jN��j�@p�rE�}�E�.؝�sO?S̎�$cBb��M!�=�̓q`��F�_�-��	���A�T����p�Xꒊ׾~�i�p�İE~����5��ez��F��k���^n+��L�m�{��M�Sy}�*$�z�^��h`z�b�F,��n���85xօ'���ݳd���&���)�d㡾����G�s�L�� ?��5��q�܇��
����RE�uc��݃'B��o���:?3��H:B�C�.z�Ի2�XH��6B�g�t �&��}Ei^}�Cj,v��ls#k�;��FV}�]�t/�?h����q� �͠6^�<�w�Kb�4h(X��xX�B!z�E���b�=�� &ߟ^��4_B&{�m�JR�S_3E�k�8
|a�H���EFԸ{�@?rw����xT9��-cb�:5�m4V�o�C��|���U���4Oq�<	�v0�Q��!;���Q&{A�p=����k���z~>f�#�T��IK\�;g9����S�y2��7�:_��\Ä�f�D>L[i*�5n
Q*6���LϽ�w��[� ��ӄ\E����IM[�M;#<��s9�u$&c[d]w54�W��Z&~aa܃�?���%3�rh�.��t	*D	w��N8�%�0�f��3��@sΝ��{AZ$��(q\�ꌶ��9��o�}M`_R=���'e��K���;������-�Ў<!��nQ�����#.��Y��|��''7����4NW�Ǯ5_~�'�rY�<�8"ð*��&E�YƄ"���Ԏ֡�r*
Ġi��0�k���~����U���I8�J�i3;�v	�y��l��#�Tٱ}p(������H�N+OT}�g��o�-����ҵYH/����s�I��v�y�aHZ%glw���?��s6��w�KoY�C"T�N�X"�DM*ݲ��v.mr�S�9�3p���F����?I��#p�a(E��v�#�� ��F�F���+)P�'�C�]%)��]����:����J���E�N��sz:�2�l%OGB�������@����sJ�$��0	߆�m��6�	a<�Bg�C��v�J���пza�(}��"���:$ϲ��v�m+�,�Vk����TA��*��q�N���=�s�8� ��$��o��Lj2(TE�c�1��F$̌V�%h��/��eI� ~q��uD�V`����n�8�m]�U�GnL�W@rW���sq;0����\U͵�En��Lgg3���g`�?(j����GJV�� �U4Vy���[�y��f_q�ւv@i�0��|Iߕ}s�zd������_�獪�;�\v�o��	~F ���bem:�pq�n��f?x
�(��C\� Yhj����7�h��dN��ʮ�l��u����p����(		�9�Я5g��=z�r��w���v��TG���d���
e>�x�n���ai�YF
&R����x�X�V�.�������+HZg��cAۆ��|W�.������  LH��8���5����j4��U�q�ߑZ��*��05��wJ�H�T!G^��Qz�~�<�R�CU�;!��v��#6��pЗ�P/(N�rC�Oa��YM$����rE1��^1�+����.<��#X���lB˝�`F�C���H ����g�)�|�o���̺#��}���^t/xu,���w+=�P��>��cV�ͮ\�D��	$-e+�k��T<VW����Z��Cq��Β)�2�~0	l����A�4��R��f?Ë+:�8��ԕ5��i����Xb}���Մ	��.N-V��2*�T�kK5�_oB�USd���=�W>Z�srN��:�#5ڋ87�* �ANzd��x@@��1�`:صl��;01��OTI����& X}d��y��+�z��/�G¤3��k9�9�4И�f���ʿ�b���c�J�~l*�)��9�/&K	�M����%���u���[D�6�	N8�4�qLV�H�SPj�9�.4�_��O͏t�p\k��u�R�m{�X ����@Q��9�����ٹ=��4îXs�Q���_װ�08��F��-���=�|���-|�f~풲`�m'>鿛
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n��=Q�8tV%d��L!v<m	Hn|�������!w�N�Fb�o�F<*Oe����1UR���j.����t�$�㮟�%�[$ ⳟA��Sl�R]�6�芫��h]x���wvb��=`��:FB
�d�U:���|�T~�|+,�D���^��nt�7\�
&������p�m�u��q��7�v;��kt7�>���b��VC�3��k���`��X~7v��؄��	���Һ%R��;�'�����x���Y�yg���%�F*�R��0���| P��I�/!V�@�9� �>Q����#	[�42�f�Kח�Sg���*��L�i�4�N�y��|���!���t�IQ�H����'헸�$;�����k�L���N{X���A��u-1����O~7]��)+2���Hĩ�w�:j?�"�S�jt?�P�P���J�<,HI8�Fӳ��w�;$e�m�M[Q��Q0�N/PŻP�&+���ș��E>�B��[4�b��� Ga�A�,g2�4ڠ:Sx�N^_zSs/���M�R�#%<���?�G�� 1u=C��]��܉izG`*|��!�ѭ��Da=�Z�J���1�*`�unO�+0&6`p{"7���p���Oh�����'����@M�����popo���9A�WK�7G�-�4(/br0D|ux�S�e;"M�ˮ����K����M�
?'_�i�jC	�8�Mg��/�y}v!��牱?C�~�	�_KV��_o�ΞjP�q�9�p�[�q���T��̈́���<3T�
�u���|�zB���xr,����~�uY��@&ws����X�����tC��ҩ/��E��8�N�@|`6�#��.ƌ���ߖ���q��>���_��9"�˪t͝n��ي��č�n�e�E�q��i ��Z�qT�&�:�U��԰ �u�5�
���[��"����2�j4���uEc�����΃b�C�R�;�:�$�AS%,\D�t��Pn{?������v����m�q���:J�o��
�ʘ�����z��6��mx#ȀAxP(��j�g�SZ�W�tj��'qׁ�6�����n�$����7�Zw�6��1&��A���{޽ʞ���Ｚ�!N+���:fb�r�"[w���?��͟n4�ŝt��Vk��+x3��N|1�O{E����W�6���z�[Ә�p,�z,��z�iI�g�}[��<��q�|�^�M�����V�_�oĭ�%PI*�.(����C��F���r{<m�NC@����B�E�k�V��-t�{Xm�[��.�g���ɖp���mGAqF���o��e��}��˅Kl�1{��t�����<��}����NLd�]������\��cҐt��e�y���,�~C8\��(W�.��G3������9H��,�|[!������:M�s��r(7J�]V�P1׊>
]��г��?�k����VC�����#�|���/�=KuF �i<l���k?´���HG����e�<��˨��l���`�z}�88���Ksљ�������D�|8�����qQ0�<#�vJ"s�ԑP�����&4`���hj���)��w#��Dqu�1Z`m��|Z���%���cK���	3�-��M�j�e� @�_����"���v;������8N�#�}�赧t�3�a�i�/���,X �G�6���=9��V�F���������M�z�_k
��|�ӧQxy���<)�-�q�.�_�뻣�8���A�&Q�Vb��-� ��|]����>��L�xԝ,����r�)$�+�n�}��j��?P]�(=5V�m��'��]+Y]�j��FGbs�
[����"N������X��g�`�������K13:�>;��5�+�ڜ|�r���.���h��B�\���ld�'O%���[]��y�8�O[�^e��$��%XJݞ�N-h�cj=7�M�Ɲ;�ϩ���M?���֝(����RB��Iܨ��nS�V)��"2"�Jd8*M���=]���$Fg9�	#�`D9M�'�-\��i��&��<��	��%_5o�X/�/��T�3��|T������Щ�C�#'��1�T�ٔ�/���W�w��%����O���ѫ+ �~4�u�uiLݘG�{2�J	�1�u�/C��0	���l��'��hK�Z7X��'��\fvT�����e~^�£�ա����
H����(y���l�J���v|������b�"����?@�נ��8��4�	?�W�t�D�%F6��0�?n�#����\hf���<��YY CS˶̉S�24mA�� �t���F2Un���Oբ�(��k*/�����x��p�_����
�GE�����3�����#RI቏��x�|WK��:;g������x�YX"n����+n&��uB�m��8�R
�6t׮�)����	(9�W��m}��.�����Ji�o�o���R��8�E�+�#�s������UQ-n�Fǜ�ޟ�����E�i*k�{is��4.�l�Uk�p{��nk��Z��N�0]�W^���u��gf�M�y�]��0�����#������k�JDl�M�?�(���!5���2.EWV�*�m0>��z��)�t��I�˿�$��U���p�|U�����f�5`9T-�H���l����.f`��� �օu"7��#�#w�a[(��S�Jp��b��c:���%q����d�e-܉7����S��(��#EEt?����l�Y�D�q	�
���y���-2��NA<�"�|h���]�nHkvZ��h�1��U'�vziʧ�[�& ��M;Tc���vIg�B�v�H�:po=��w+0�z�h��]V�����.U=��\������Q�Q��T	��!���<�ڐ�����{$%|q���eq����>eN�����v,g�G1�g��r6A$q�"2�w�+�juZ�ٽ���N4:&j�C�-�lJ/Qmf҅�g�1��[�̾�����h
;e����@��p�a����:Nk���&4���"�
eC��w�1"�����1<�f^u���T�����S)y���W��z����
ɳ�<�ˌ�ݬa��$2��������_В����.E4�/�4'�0�aD �*�N�a��>�iI��t�M���{�?c7(	=��HgE�����Z�
���K(ik��_v���^����V��-�؋���|�������a�o�j[��z��X���ZΚ�����r�iQL�S�IT�m�w���O���_c��V�w"���Q��F���k4ۇ���������zB,�E��!�5.�3�k/�ݫ�g$YQF&3�G�>d�Hilyb�9]N�7͟��ю)��e*�=*����.,���]�����(x��W�+V�0�o����h%�QOY��4�U��tdl���|�`�l���P�
���r�lG X���Z��0x�!9�P���I"����<ԣ����tZ��r�i��Cx����J=c��7n���c8f媤���m)�9��v�aW��P[�����7�\Ƽ>�G���j���)��a�j�\�_b�(���30��X����F�����C��?
���U�@gѨ�jN8*Z�c7�]��ߖ�[A<R�!��{iڛ�p��V�Mt��ܹ�!�ې^F`�t��7(d8a�P=�{���_�ס��;�픑��ܶ����~#k&on_��'7V�����{�0vhɪʈ�謗���PW��/����G��`7ʹ����&^�9�"���6#]x�u>R���lK)���$膓�/d&���8�I��;c�C.�j��d�a�����t�=�I�d��z7r;�Xv}�N��f;�.K,Ԫ;�!�.�I�� �4��9&�(��sg���~ɭ��	��&kѬ�Q�����g�̌gw�KS���JX��g>��D����U��^�9Z��o.t�Z���7G� ��m.!7牣��SyPſ��%��exY���]q��=����4�7��_'_�v7�|W����R�n3��6Q��B{:�a����7���.v���3yu�{g>�k��ԡ����(�A���Q��Q�hm����$D
��L��]�����L!�Of��t�K�BU.�x�U�%3r��,�v��T�e�x���m��}^��F"��0}�/}c���]�ʨȸ���%����n�i�:�������q�Y{K��TP�%��?��,|�[qzO(��p9�	l'�yA�Hw��ۭ7C�䫣1��WA�'�|6��ݐr�8\?�Z�񉩊���Ѽ�/89�
����TӛC�4N��?	��fr'�!AĊ4�="���cjm� S�B��Re��"SP�Vǚ�&���_T�ŅD˴Xư̓=�9��O�(�>Q�T>��5�)�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�
#�i�MS��Q�
<B
�t?{�^�z����$�����Yp�Z	��O@�/iO۸�3�����p�`��#���+�B�&��Tf�O�}�li��x������2��c$����<Ԡ'��Hb&�[�q8غAC
f������8��]vʝu����@���-@�0{o>����;��9���1!(�g���?�
C9
e�Y�[� y���Ts���b��Qu
�;τMk9'i�=���h���\='��c��+����墍�n:<��UN0��k��<j�[�ȋ#+a�ݨ���Y�z�cc�PK�2��Cz�]i�5�:��Z�B2��w�g���A�ynp'��Ѻ~��{�F�XQ���$x@�Ҏ�����S�������@�*����Y9��R�f��o��My�=�Q*�	C��5������1�hG�Bp[�9�#s(�8�6F6z"�st�4�r�N'��"%qj?ևZ�C�
Y%5E�:�mB.V�7�P���	��j�.�7o�^�+���?U�5������ 9f��b}�&��AOQ�1bn+	#��j����)�oC��B*�
~�+Q	��SE��[�!���h�v�ʇ�g(�^"�� ^�|}_�B!��j0;1���|����POV�
8:�9K���U��i��nn��%2�Ť}�Z*ǵ>ˍ�	;�:3��O>������?�.'�=��
C�Y�*k�ש��LU�d2̇Ӆ�痡H���װ2��hE��ā͆"2a~d�l0�ҬD7�2����L4`5��������d�)���7B
��hf���܆R��P�p�&gb���guvo��X9����wEFɭJ�_�<��!8���?	���W{t��e��=�BJD��+[��Ĩ	�Ult^�ڇ�7�|�
E7��W��0�f���=	��� ��h��8��kDy���}Y��D��Ħ¹ތP�)�j�ş$D�����"�n�|���~�bc���9���>S�)��������^�&�h�� �y��"l��SALX� p'����^����$��%������bGl6�Y����n��r��r�?ܵ1�?��ڒw��h�w4���5*����Qg�)�ok�Ju4 ��,�O�Շ[O$D�x#b;:f��sD-�*�j���p�7s�/hť������4˰t^�Ǌ�SJ��}b�Q_�j��*�FG�����'R�ψ�*������
k�P@NUp/Sqf���5�V!}=��ū���?��u
��H)��-��բlX @[��g�BYۍ��2ٺA��dnR��r���
�<�Ҭ���L��4 ��HB��L���͜}��d��k���3���q���� X0�%�RK�p�"_��	�����lJ~��%�c���ֱN��~ �H����~[�Jd��6>�|��%[�F�׶��umN1�r ���&������k��:v$g�Pų���pt�� ��.դE�B����$�U�e[E�r۬t���Αz�Z�{�� ���|��+`�G�!��h��9���h d�<�iQ�	�;T�wȔv9�C��9�p��bor%���>Q5]��|k��_���<�8V�¡���^�`��4ՙ,L@h_ ���f����t��n]�R���)�	̛��Z���΃�C��?��2����l%�\�_3�ćwث�^q��T2��^������]W����B1�6mYY�JВ.RX5r�F���: 4b�1:�!.��M��zD��!'e�w��4^=.���t��b�e�7��=?���:���-�_��=�~�dR�����"�q�V^���a��s���+,1k�VzJ��^���0U��0��}�܏Sr' m^A�,B��XT4q��@g����)>�>H>E�u@��J=���ٚ6��xN8)��yv/��Ya�1�櫧t��མ�SSH�������F�'g/�Z������Z�Y/{J�����%�M�a�z��|�d��[(Wڹ�J�Zς����S8){�N�5�3������.��B���匃k�����H?���[�P�j)�WeԮO@N�t ��7��������� `H��B9�P�]���^t����̓��kkhy�u�P$l�: 4 �z����|�<���������	?�T������^�C�<�V�>�f55����y)����ڳj�\��x���>� ���s�FL��j!o�m������9y&�7	
�I)l@��1G>p�S}�`V�F>:�va�N8���6�}��&r���3B]7Ta�!�9� @h��5�&��� �����=�wRC�Q�>�9"�Y)�\��߽z���&����uJh�b����O	��v�"�g� ��Ђ��EZ�x�5��dPuüI˖�̡�_������O�3�B�RX�4{w��$lg钂S�N��n������	�G�yЗ�K�s����_�p���r\tT�2V�Ń��d0�g	)p��=���r�5Pw�4��!���೬o�����q��Obcq_��;�^�	�h�� r�f�r��"U�dz��Y�Q :'��uX_�A	�)69)����PJ�Z.<�ec�M�j3�B��R ��RE�cø`0���A<���+8����&9d��t^e�����
o�2M�*�=��ϴ��h;w3O�F~3u�\p!:��O������<��o����� N�_�/Z�x���m6��#;�UE2���T�ß"���㮕Y1Vj|u��[k��I��Za�|N>�II�;���?��X��:S.N��,4�q�+Vk���zb�ĬU*t��i��-���Oa�l�Q/���|���\�flYg��: ; Io���N���k�)9]AxraƲ`�3��Es�0�=���#��{��V�ƿ)�/�̩�O2	P�7>��V�I�`�<a��%þ���Z>�z2k3X*��RS>=~C�F�H� "�>&���W�6����������nm�V�kamg�$Kw����ޏf�p�n��zю�oJ�g0�o��Z�$^e��.8�4�@��褀��"�M��I���ˆ�����Z�����U�U�b��Y�BH���\v�/�����U@{I9~�9S�>�P��'x	�b�0i�by���^&��S�`�d�-Q�-F�j���d��\Q�wK%;B�da�\<d����V�ڎ�C��ۙ����muQ9h/O�6��璡���1|��ޭ��V�Z��d|*�I�s#"6Hmo9a �3 ����<��`��_�T ���G�����6��[C�G4�Wļ�����u�,|3�_�n����}~q���Z��"�
:�+�%�E�+qѨ��iB�C��E����]�,І�����8]CZh��@�?LC9�Mcɾ�K'Z5_4�����>n��DyJ�%��a'�j�����`y�X�������
]�ي6<_�8�z�2raZ�O�=�9��)&
O�Φ�����J*��e�3D~�Z���B}qi�q�F[CP�B��c4��$R�	l�2�Zu�e�x�T�]6�@�M��Fפwƨ�m�^<+���#D�a��c>���GLh@�f�,�$Z	�� ���8ﵻʁ�n�k���mĘ�����m�X���]IZ�Cb���s�3ds-�[���9����M��%��3p�FV�[�Mb������U�8����s7�|̖�u�|�]���j\0�W]hH>�qw�w��}CW�~�IN6�LQ.;�Ui!.��j�(��XАBp8�ɥۋiۖ��~߲��2�>8OJ��n���Rߪ/J7�>�*nͺ�}��������Py����x	>mH�Eb��wbp��v�b
����������p6cc\C)��r��{K�Ǻ�〱��߼��X癓��J���o�l`bID�`��^B �5:Ö�}�QȾ�2���5�D\g�C���1	Ë�(܂�|�z�=�oX��q	,
^�ds3Tg�X�w5��L�h���x�q����P۠ӿT��y�S&l��|8pbI�/�^�1>u	cT����x���VZ|"x�&�9�%�-Y{������姗�;�ܖ�~b#@��Tv�5���<��93_�3��C�4.�*���S?�R�?tW��b~G�>�6���*�L;�$��U���5�RV�R�ݣztB�����o6c:�	.X�
���]�`����"�:T��DP4�<>���^L�E��+7�Ҭk�=6Â�.��9P��i"B�i����W:�eB%���&��%��=u���鸮�D˥��_��ބ��� �rU.}l��d]0D8PV�}���F/zl�,�X�9-cD��#4��{3 4�r䟃h�/�6*/�t*8�]W�?��f8BU�K�F����]��y;س��]�=p�q�� /Y�Hy�*n$pjC�����f8��I�X�S�~��M��+A�V�K�MF��f,�s3T��������QY������G^MA��AѾ���HL����q��Q�9��荝eF\u^�����HK����I�ʻP~�l�3��)]~=�Z�eJ� 6W3��R��q�m�Ea*�Lȯ1��X���<q�?9��]�ͦ���C��b!~�Z�L��脜��%~:-�ǁ*쾫���{8�Y�\%� ��QT[��� OY���9w;�1���q��ӟ�^B�UX��IR��0.�y��'�饏鑼:h_�²����7���yw�!y��T�o+5BKH� )���1��A}�۳�\d�#\N9��x�A��lI��F�2p�+���jB��<�HbZ\�ᛥutc���H*I=
�Pr�E���z{��:`��ϔMIM��s��1�M����~�����l��ye�'vhǸ�=B�X��'yz�Tթ�U�YG�:�Y���`���y����@t�pe1�����{t������a5)�h�*f�`ze����b읺.��q"�yy[���P�c�+tkS\�R���J}+J���(�mS�ۄ�@_νb(E��5�x�M=B��vF���(�!�bJz���K�e!���G'�-�m3)���r��6��I�iy�ܟ�1���^�"/��Q�+�3`~��8���~MoD)�pD��#��Ɏ走�ݛDۨ�F�6�S��[��mO����±0���E�6`;Xvj�h�%=�~T~����Vh��.l�tZ�d%�A=[=�ݬ��xƂ�7����3/�\��ayƼ�U'��%����l�;����B����m�p^�����h��ʹZ�qG�l��<��A�˘@�ʏ[���i�:�Ĭ9���g��^��	sD��v��x�:;_�<~�,7�DV\e�e!n�!#���,�]M��fA%�Y��?v��pb���ϔ^1�O��g�}*mp�z~��� �̈́�~W|@���Z5?t�:0FO}Y����0��X��$�&?̎��W��2��"�b,7��{��a���{¥�V=��=z"&�@MZ�jg����Ș��G��	R�6,�}������̿%Ӛ�I�WE%>�k��߃�Vx���o��90l
W9��d�� �b�	�ϓ�w'�;] 	�0���S��D�wi���HP�ʔGo�.�~n\��� eE��W�J,�f`�ڬ��G�
S�£a_�6��7���t�BC�C��s1��!�'V+ra�	����/��%MC��}�����pʉ<�
T>�V��L���O�2��|����R�ώ�27��3��ľ�N��6$����H�oԀ��(x����|���<���4���~��C�C�N��V�ϸ�O���߈g@P���J�>5�����]���OأR@�x�O���q��=8?�p���!�~ �B$�VP0�����B2��D�ϸ*�j��9&*��)�0��� P(�7V3�f(z�t��y�w4�˺���ݗ��Pd/�}9���z*��q�+�5ζC�^vI�}#��?��.�KҼfતAg��Aa3'���W� �0�-��}+aV�)�8�ߍ��R��_�B9���>�/z�}�Ϸ��AGӁ"��;mC����U�P�vGi�LF��je�iA��ʸ�x���IuguWS���m��]�+t���qK��=Od!�D�h�����w������ 숆 �g����&���x�0��w߹"[�>���YD(���ſQ�*DYf��M)�o���i�`i�i3�e}��]���Mʷ�-l^����]#x�ۥ&O2���������6�����	�<H�����f���F�L�Zh{ii^l�7H:�y�<�v�b&����/!��0�.��)Z���+�Q[?wh���L�m�
D��;B=?���JB�z*hƑ-"�E����A^��aQ���@`�*�����y�2�_[�M�'@�6-��ڂr����'��k�ZW]	���菲M�C�|�eg�vb�4z�x)Nb5�[�;�s�����շ�&py�%��k��l㽳
U�
���E�ߊgj)����:M,'�Y�Eхj����Ô�T&���"�L7nMJ�N0U�=y��7W�r�f��� �D��L��;��?����;H����F���r��X�q�+�/��@q�{L:�#�.��KK��擓�Ȁ*:�/3��^/Y��t�{D	T�$D��7㚒��gg�2�a�k4,��G:�6�xN���c��e��:@�Yܮ�1m�f�-s�;���z[Ew�ey3��\'c.��/6O)�[g��C��4��I?��;��V�ŷްS�;��?<%-��$cG���Q����o'��ɴ>��[�UCPq�l�N�Ӷ�1,�0ή��no��s���*c�6! �ty3�2�}]�쵕G􅿆�z#�D�ܪvb4I�ͧ�(�:��V��>���x��]�^i孼q�(b�H���(��<�,N�	�V���A�H�������ٖ� ���|�ܲw�k�@�z��ss�K�^~�h�jC%����o�(��ӏ�3^���˦��:�v����~�&���l��)�f�}��RM%O3��~s.�F����{��%:a���&!��l��<�>�)��B��g
ϊ<�w�����/3���k��Y�x��	<I�1$Ht��A���1=4>C�F�}�FL�ň���k��'���F�_�%W���4ܤ�
0�օ��T�?�@�t�8���T`P�dF�>�x8g�E�=�b�@�Iobl+���M���� *x���Ӽ��8�_�ҨfF_'����N��p#���髏�-s�p��G��*�`C�o� C_Q8�$5o��`6�1Uݓ2���:��#'R�w<�R�C7Ŗ��5��Es60yR}$�Ma���]9�3qڨ���4g�/Ba_,}	�@�(�h�Ѵ�굄���G��n��7 �����$z�A�#Ɠ����39�IC�|n �pI��΁=��R�%�����
o��)���1�𡧨�s��u�ıoͼ��yRf? tJ�|
Y�������CD<2����A�~��)D_�w��[�Oż����Ò� L��� I�*�3��PUh�ưN���d�5���g/�Wm{e��i3M9 ĩg�,!
6����6m����k��B���2�=�)�Ĺv��{��媗	H��v����£O?�O�"��J1�	Ƚn\OQ䙲�k�$�U��7��tzsr��9�8���3$܄8p:\��b!��]/Xɋ�X4�g��y�h{�*�o�IϺ�vs�!{����C�.�5� 7CG%�P�G��
G�s=5���V�!o�Ŗ\6��L�?����ܾ�f�o(=�F�:�
Vz�n�T��؈!,����Z��,F�fSkd�	�.��:�@��w��8ʀq�6%"��Rܪ��5���k
%����XۨN�V~m)e1�w�O�s7��`��_!K-Ϙ�m.���?�d"GC�e%�1�ƥ2E*Mٲ�k��W�ӎ��?g�٫$s?�}�����Y0C[�\�h��(tYT-��x9��y�>�o���O{#����͚������ �K'GH��ڳc�L��I�)���d�s�'�:G����wx|(i�vP����@*pT�U�ޕE���xk���b�Fl8e�d�ŏ��Pd�Gٍ=)oY'�\h���;6��m*J.@i�����<�#��$��w�� m��;�!��<����b��l��vo�r�t�/�/S߱��(N���E��7��
��������A�m\������ooWx�����`;���vF q%���9^���ߝő���!�c��ˁ,��5%�O����cQj��ݿ�4����[Q�")���~#��ɔ�+�����q�[��Æ��DY�n���׌p�*��<<�5��9����Ra��a��z�8]BgχN~NW��Z���vj��/,��G��St�
���*G���4>�5}O�fB9MY�y��<p��se��l�]��{��0��Cmi~�H��|��9�f[R��X�!���
�h����0��|�d�jq�G��#QQ.gYK����	�}뷺{g�I��Gd��#��W��k�y
��z		������zUw�	n��v�uFD�zX8v���O!yp-�x��Nq���s`�I�%���1Vd�v�j+D�%մ��L�|��`b�(�Hi��̃	��:Q�p� !���I:Yd_�eSI�1]�M�;b�\A�]���I&Yq"�v֬l�T����$w�[B&�(=��e��\��/����Ty�˼=��-S��5�����j�(Z֍�(����c��	�����y�I]Po�N6���{X�Z�f�������B��un<`Zr�>�a�T�.�7�KdZ�R���n�&�t[��Ü�5�% �輪B��q���Pt�&�D�JVK�RPN�F�X���nm�}lR�5Y<�0�g��j��f+�
�d��$+��c�Xd[LI)�o��ZȻ֥�eу�= ��`#���3���4y�L�+F���ZHor�����>=�s��
'���	AcQ�mf�։��Cp^9���*��)���I��J���L	w���]j)��'���G�7��
��dKrgGV��MR�|L����͋pC5�{>��`�H�\IL�#�	����E��	K�S�S �*"���#�Ϯ�9�&`�XRΫΚ�E���^���P�}7�!�J"�&=b�?L���|.��|��pQ[�6�q�׆h�v�QٔB���?�/w��nsoM�o���5@��O�o' �8^�cD�S�go����F
0��[�u�F�5�vp��F$5�7��-��S�	��nK6��t]�2-����&�}�lK� 3�C-Ӄ��k�q�x?ۘ���._��TkZڍW�P����x���/2h�p��?�'���oB���M�ݢOֻ��̮ɒ�X$�}�ui��IG�T�LA�p�CK4�z,��}I���?ٙ�a������i�ue��Y���3F��%JZGd�CƵU"��D����y^=�cMy�����C'F��$ؼ��&�jۧ�o��Q��u���>G�+9!�L.,��$U�`�}r�oG�G���h�%��.S���#�j��9���q�x����.���N�09G6�� я�v�߻�U��`5�4>se�_��@`��.��'4��S�kH��ከ�u���Ϗ�Lu,�!|�c�d.����B�|Y|69����B����2�q'm�3��ƴz��j.*;1�u�;���(��_�K���y)��e��J��[�:�D�۹(;�f`~���(V���N����Z2�:ƼƬ�3$8�"�L!2���3|��5˧��Kkz�lY7Yv���s�[����гYa��I�"�����ه��x����$U�B�F�ͭ�,���a"�_U���Xa��v�;��/�X���n���~	���`�ɬ���he[�{<��6e$EV�o k����*��-�>'��mΨQe����r���`�n�PO1�!ֲ�3>f�H��	�A���#~�$@*i��I�@�f9�K"mvq:z=�%=_<�>����W9M��n�5�v���D��DH?���d�fi3<	�^�,w�ҁ҈��WZ���겶��-�20�N�R�
ڍ\&��{�\��P�C�.is���WIY�W�zD��k�������"[���Φ�R�q ��ݦ��1�L���g�C����uu�&+����X-x��5,KC�>4{It��I�u䤄~{�]ĆR�\��k���ȋ�<�}=nՌ�� ����m��w�y)���Ѡ!_�<��?��W?ˡ4AK��[8���� �-o��q�k|.���%��m
�?� ~����21i����M��|P薚A�]:~"�^�k�N`d���EB�&"��J�NWo�>��� �W�-p-� ��ňr��úF�����Dx�(�_T���10	/�)�U6L�9��D�������c
2��^�r֨���s����ir�z���������6Y���ua*�p�EMe`��urΑ��D�((�^`w��y�%E\d�#;�p���s�g3�����d'xm�;,��	M#:ݔ��RP���q���˗�q m�m�=��9�O��8���_���}��T`����󩇰�c��Dy3Z2lO[=:wK~
��-G�n�4Т�M���!�Nm������0���ye���BݠN����7����u�d�jr��K�v_�WWx�(��O�_�穙��Y����f�ʺ}'_
�(B�Ɩp�'ԗl��K�3��ʆ��^�M@O'W�{����v2zX���}l��
����A��eO�W���Gb�5מ6�r�p��g�qOӌ\=����A>衐%�I�x��:�~����k���n�ZQ�	f��In��{����3�P������9ko�Dj�^W�.�菼P�?���x];�9n���\G1����Y�K�?�ƥ��S����Q��|�(����&N0����R`���i%�x�����jCt�3��q ����u�7ϓ;��x?o#T����V�K����pM�c_!�p#��E� 2���1#\Z)���:M4ʨ�Q�����	�&' co��sf�����iBN����R���ad�	I�����V��N�6������ө|f�l��;�	�4̙E�g�o�i��c�� =m� 9��r�Z�D�В�J�kS0cQ�4��W琒zͥ��A��vS5̥WC�p?c���{�f����}�b�H��ײ��#�}�J;��h���}�#��9�y1�8�b�i���O �p�#���:�J��P�0���P�v#���U�1��2f���rG��գ��;Ř݅�+����k�\聕�[�����|���@j�g����ʼV$�d<H�m=4��vN�+y��8��*ZjB��i*���a�HS[9Z1 ��.���.K��J�>F�A����l$���:܊H>D�?U�m��7�t���*ʊ0�/����>�GS�{샯�Zӄ�j�#���`�g�ipJ���v�;L ����X��4��],Ҩږ��b���`1k�����p�d��t��1�Z���p�u�C�:r���D~�*��o�����~���%W��aӡk�s�B��ܔ����A7a���ܾ��q��\�0����V�s}�bxq�������u}�؛re�k�L�<�PPQX�^��{}��ԩ�(I��zrN��PJ��-����ؽ�p)��,�f����5���?3�}J7���\�0њ�
N�k�ٳ��JӋ;�~(wy�:=�<$���A6	nW1�/rQG�OP![��Z׈���=?��$r�Jb�]A�N�o�m�\\�A,�������W�7���o�(����d^��6��}ӡ���m�b�T�{忺�/1�������D��ab�� �o��:.���=k	Y;�@��!����9����4�%�f�Ĳe^J��*ݙs�ECk�H<Y�{��6Ӛ�Yo\�@�v95]\nS��M���Z�t­�j�⩀�|�5��̠�E�h%�v�i��۴��}:%�i�av�@�y�Ҙ	���0-/c�gb���~���pdpj�ʎ[�Wr\N�:c,\�N9�p�SC-�ǡ���@bE眈��˪'�<�#�Cq�<�>�h���#�<e�����a���Y�2 I_T���U>y��'ܨdնU"�5״w��Hٽ2�k�>��k]y��[#ӎq!Q�3�a*���%-��!�~Z�)�}8c�j��T!�;q�M@3��K�]`cy�b�,~����9���qFw
��Bpu�kn����;�(4~v#͹`+�*�R��ײh@�cY�rݏ.�l��8,��)i��e�K��v����c8z����~M�M>o����@�Վ@����m`���
�m�l!`l���sң=�2��g�*��{�.#�	'c��-O�Xa2��_jP�:��m�eI��RbU2��1v�}/�25�}J�>d&�}��@�"�����t5G���	�k�b����hv���>a,Y��7�ls�i�t5�:�JO'"�V�1���I�s��z2)�T����G��C�:���%��P�s#���5g� �s0E%p�{4}��85˝ʫ�*������gmd��Ü�������j��s�:;u5!����P�v�Tnf녣���=�6d��i�Jz��|�z�3͂R1��f~���Vل���`�9���b���P~,o���n�um/|����_}�)~V�E2�g߹ 5H�v�JƄD ��/���0˧j��r�%�5UWSo��9��r� �A��rH��|SS�ѭ3H{���<�n�]��Q�~l(�)�P�gn-qW����Fp�B{�� �C*��(�\VZm���b?��ȡ�R
"Dxs)N� )A�w�ށ9x�n�&�1�	e8$���hH��$�i�<�1���ɞE�<a	��BB'{�yS�Mڛ�Z 	��V����j�"�{�x�F��H�G*~m�6Ռx�J���ֿ_���9�6�fՆ���ؗp~;�Հ�x��u�e�&��r�Q>��٥5�݀TP�+ǽUϔs~K=��	^$�DR&Y�%�'�.�$��p�V���V���ď�|	�ǱK~Api�<����?Y�t�~�ǃ��'����K�f�ht0���Q.����/���O����1�#��lm(6*�a*|&���=���Wd��9�=u)���QO�$�ӶL����b���_�E�4����t�В�����!�18��ZY@X��کL�"��LZ��$E* �K�Jw���d- ;�F�[
9F�����lz�1���PO�W>S�hf�X~���'�)�$��YX`\�6�E��C�5��d�U=��]������O�P9��\�j��0�5J ~P.M��o��>"��M�U��G8�f�Vƌ�g�8�D�[��r��l��������a����iw�-IU`lP����O0do޶<�^�{ya`6ɧ&c"�R��I5�R'u�0�$h ��p=�������+��p����h���d�Uֻ��������F'\��7���^�İnq�܀��Ōg�D�T�ݒ�>;g��p%���d�:K�;g�A��6�(��8�}��D	�L�g3a�X�nV��q鈖� �?G�\�U�(�x�o}���-rۇ�YS�7.�rzYڊn���>����y � 2����/�j_#�4�`�Ω�� T8|�-��|��KRR�S��Vyz����(6U�tb.q&��U����]�h������D���<�.��#/�s�����H@F�֖�����SR|)Z(O$w�Oghm*��:��u��wB�}�/���0��<�5�z]*_r�rPߊ�w);���?�{M<ɒ��g�VV�<�[8�SAgӳU֤S�ʆ����߁r�'��=�f�q�v��,��_2�O��H�HgNB X|�K�UѸi��/���q���or��\���Gע�����x8�_pJ�A;��ӕ���(S�:_��7n�;&�5:���K�z+�����׽Xc��ioP/��\]��M�z<W��7Gj��Kc�߼�/�Іq`�խ�j�G�n���>��_"�}����\V�X��{��Y��#C#���hS����}�S��.�i��H��b�T�d[�j=||��A�?41l�-�6��
�y/m��5~|J��?已�wP�B���y�ʵZ��+�j���;��!bf;-��|�Qô5�7s3{���z��������v��Fס����Lg���M7��}�	Z!I��W�Ʀ!��'<��_nҧtn�Ш�������/V��	�|O��ܼYzN�Z�,{�#��Dm�k�}h@�7�T�HƂ�������ѷ�2�n����<
a���'�'8b�p��Q|ϣ}���R�_"����d�7��/x��$�,�����X��9r�W�rKӯ����LG�6�D����Xڠ:{�6 �ښ�V���DD?�Ck@P�>w�1�p��/8��8(JXRPu��k�_��P�r���k�V�qQsF��0
>��b�L9^�D���]�G�yb�S \�,�w�R�h�R��#�B�x�L:�3��韕�� .����|�?,��9�hu6ny{e�/�6�����w�����J�k4$�X�{�k���sp��/3�Ff�r7�Y��h�ra�� qC�Ϗ�?g�����'����&|s�IT�W^���/�	fq4c-^V̍wJf�|�SC��ͩ�c���7P�ϗTT��>�E��Z}Ӭvop=�bZ�z����Vg�#
�/��-rMp"��){�MN��`��g7��!<6")��,��@A����G��"Ʒ' �(X��yB߀�7���,�GLe��i�ַX����}�5r�(���>v4��S��!��L�!�,'5��\Mٓ��~�y���D8�e��[7�<)v����lD���֥om��ۃ4�-�[���E&�
&V�G9�)�����3@�Pq ���R�$]?g�1g�i���.a��C�
���`c�x���q�@~�A�_$��qx_���vƀ�i�����u\|�5�qЗLU�#�p$�v�������3�UyjbggnBNB��q��:L�f��+��p���p;O$��h�;Ds'O~d���g'm*&m#VT]=�tF?��rEK�~����'�H��,��k|i&�{�>,5���|حԈ][�:���Kx=XCς�S]WQ�ޅ���yg�%$I�ip��%�׊����-6X��o``@�s���+��T�,��"R��)Z�t%�b�����'K!-�=U�|�kF���!m��%����I��x��Ո�0!Udd�-J�ȹυ��{y#��P�.�=4F��͖�VY�|�P �ҵ�^8��!7���� Z�~UqD�A�ݱ�$U٪q0�e����5�$�L�L�6�^d��M-i��ޢ<���k�A�gL��L[6�Ȥ���*7t�f0�'�	hc�� y�fh���\0=H*�x�.j�QF����;�Έ�<��5�a!�B�:0��s�_�*�n�?K|�m��BAa>2b--b%a�k�����3k��{��b��9�᳍��H�����{r�5�*��q��w��ǀ��ڨ���>ק_�1q3��*庺�z�)��I��o�1������X}نQ�(=�������@��Β�s}��V�)\FP�-�Wm1���4�T�vCjՈ-�ˡ����b�*]At�O:t%�v��oN�{�5�m��j��4�����K
�J`.�)|/n�Mm���~������Z�>��m3+ض�瀉�-��jf�7p��5E3�	S�~ۀ��?�EcR������r��#/����6�:kQ�*P�Cn 0K$\5Z��J�ޏ��~�>�q8J�uT���zU��L�������p"����"#-�Qe��������Jү�L�*�&�����!�� ��o�"���>��G��"��}��7KRż.f3~Oc��DIz!�o�{����}�|�)0��f�_%�9�a��G��lf� >G�D���hX�Ło��_�"~mɽRd��d7'.������M��B��>_h�.�.�����ͻ�ā����r���m��oBf�f2�n�7~�'����[d ���dX�Vٚ�劒�#iZ�D������[,K���M����f����N[���N��� $�Ȟ��!�P��j7�*�d	���C�hO�����(J���dQ5I`o.���Y��o�� �?��_�� ���ލ�}��3�jQ�� ����.e�HFk9�Μ��@<����4E�g��y���YZ�j�a��5ItӺ�N�;���\���`�P��V��}���+6�R\�C^�<�����zCEaej�<�&RӸ�v�,wT���Or���Tpk��4���K�X4mp��/�5�E�7�'��bx���D�BfI̮�r�o�F�FT�#2��n=�=����l(���,/B�>����ekr��� 	�`�����NX�t�h�K�%�!E�2	[�0�%�h��ԳRx��"��6���<@�X{rHQH�@���.�ܴ?�*JXX�O2!�=�'��.���gb[i�����)^|6DTx/��g�O��p %�v�e�6���+��x*0��4V�Y����<�3,����_=�h]	��Wv��@��dך4?Ր�_�S�(�IO�$̓�벬\�ʹG�L�BD|�L��LG]�%H�ؕ��|��l+Ձt��f�1m�!�$z%PJ�n�|?����>\�ĉ9���!��DL$�������Z�p�+�9 ���J���nD���٭D����a\�����lM�#����	�P/�Ց
��G�Iź��`C2Ts��_�H����.�<�o��7y���˞$C�.K�KI�7���Eed4@A��!{��X�5����sZ��Z�~ay�\��|��>6�t�.,춷2��@�S��#�ͬ�`�_�њ�����2���;�&�l�'����v�O	�����	W��֟�E�b%��7L�A%;'_�O�5/\�^ڕ��,J�9=���{�}=��F`<<7�U/�JVk?񟂛�6��&�����t�$|���WLyjja�4�֡"��f8/���m�$�d��~����o�2kF�?�n��KE/6kU�tF�M�S��<(U|��.���{�FM�O��ɬ���t���Kz��/���i���Ց��zE0��Y�7j96.�=E�i�{=�����V8�0�j>���e���|E�dV���V��ɪ���p�-�#��o�U��9G��J-����	�ǈ�<��&f����ĦmW�!���eKJG+@����7DZ�X�>�n�u�J����R��зgu�`�E�fǪ�i8��0���(�_�!�R�@ʥs���x��	>����կCc�S8(�X�lTA�z�*߫��LwJ�{G/a�Kd��`poyr'Ąm3��|�8]-�b0�<.vc��}�:�����=��<�����8�]P��=�g���26Ϗ� a��ה��O�8RRv�4J�����?��´s��s��s��Ne��:N�T� �l,L�z��m�rV1tWi�!�n��E�XB5�!:��� !�xz�e4���2~f^y��G�π�d��F�����>@Z+YHZ��A,���}�nM#���`M'�`�J��numc}~�&�~��Ȟ��D��� ��;Ƚ�^��W�D~z�/���g��p���l�Y��L�\a�t0����; $�u��*�$l/M������Uʰ* ��,� �.���Z�z�^��9O�D�W���&�Y��� ���4��vQ��M0�ζ��C�.l��j	�Im�RG3�~|4��Q��nF�����mх�?8������j������&䀪vSEY�#p�O�����(��r�Tkц��g1��d/�H<<���q�
��\���)D�^>��V�*b��M����BkKdA+���H�8�5ü�4�ט�$F�YS,�L�Ƶ��'9���Eؚ� �� az�E!�;�
�'vW;GwDI���
`�6�r89ҿ�
P좍BZ�zh���Y��+�$ ��~�S��+�Q�[�To�Ñ����{�-�!��(6'�z3O�ꞥa|���d�"��[鿠5����mJ���pp�eo�x_=f��6��(�OM@���.�[� �3bZܗ�R���~���S�dú1GV�c�$':�yX�O�Re�i�
��p�˄n��JCҸ(�94�$���v�a��)���L���=J\�	mfϛ��yq�7b{��c�� 聽_ö24��<�$�a���}u���z�"@�c�~%p	p�Sf��<��"~P�ҙ_�ؽN+�$�1s���/��T@�HH^��C��Q��>�+�*��m6Q��,�O�%oK�NԩAc5�����<l� >D����,��)	�\��3S?e�Z\��4E�"�j13���w��.�Zw�(؉�D��+C+Z.���yO� �z*	�N{O#B���j�x�b�Owo*/\�q�A�2������ka��? ���C�o�K�{��+�Sȧ���8Q��f`*-����=�z��<ڦ;	��1T��w1@����x��Y�DL��C��`m{�l�~Usb+�C ?�1R�l� ���f�f���1�49���B�k@��������#QA����P��	4�tߍ=�3��(!D�=�ƃ��Bw/�I��+Q:����>)	��x�44�pkS7ͅ�@����F����\�K���x�Ŗ}+����93��&�Y'꽟�i���1��L!�I��ϰ���s[W֟-��bH��I 
+�G�Mk��;�P⥡��P ��G�c�ޞ����3�n/�̇����Y�?��!�W`6w��J5@^�cN5��B�`��1x�ª��#�i�o��T;���T.	hF'�}!����Y�\�7p}�@��YA8b�f�s����Hĭ���	�6`���|��L	NX�qM�meǪF�����
�K���R��K��oG��6������;��@�+���4;O���Z�n��z���0���mO��k�H;Z�)���#�����%!�!�W�n�<z0��L��^j���t��4C��ݫP m����x�S5�7qΐ)'��E����Ս���9_J�7XN����:�RE����ϧj_\�^��
M�я���}_�����,@�pS��5�[���ʮrj Cο%�L͓&��nH	lS��*>�� ��Uy�8��L��"4B�
m8��檖����6{�Ri��1l(^쵠���mNi�`"W_�/��EQCS�|8��?غae�>��R� �|~-8,ޞL�PcC��˿��:wǈ@K�RV�ڜ��<.�t𛩳�|���.��2P�_�����������T�:NxGK�<.l����?b��z^,�$:-Eu@�*W�4��Rb���w�J	�����u��f��?⢆]GJԇ7`L���x�DK�i�%�BkJ>)���vL� ����=���;R�((�vj�B�a�� ���R�̼�|s.)��u����-�_���fӓ<�O"�����1�A�0�ӭH����ކ�+yr�L)=��"���!_U���z�(�
��5�s�=�	��TN�
;�u��iiRY0��	H�� ����ن�E�٢И9S;P9���MoZ�2DϠ����))�#�?y�X�p�0ٗo�Zd8*��p	�.B��j"�S}=TH������8����B[���o�*�Q��p����;f��e6.+����Gx;��D�tT.'e#�j3]T���,���jFQ&8�Z�楃X�/g(�E}< ;�B�.e��Ql3#��e�m';�7t���ZB|��b�I��ՔW�v�g��\��Ⱦ���M ��ڎ�ņ�E���٣[��T�)�'�S�5�_'����g��{5rZ�����ST�ع���H��u�����E��XM4�kĥm-��"��uu��� �'�A'�@^NU���(B�N��ޔ����-/9$���{v�{	P)���]fh�2���
��K�(�Y���'�>��N���v`��ֶt��yu���1�ƿr�p�§��|p�$����rKc�t}���X����>�"G�������%o�G҃;�����`NWI���/w���s2Y���G�n�'��=�E���b�5��7*�g=L~���_���s�$�+q��[�H�\���eh�+a6���J(	(#��PB��3�=9���%���r���]���g����
�:�9k����u���M������e��&T+�a�m�/& d�t�h����d�<&�4�e�$%�h�<%�����	z[z����uvT7����1`�q�!�H��Ѫ����f�	������C{Lp���-�R�O~�k�f.J6��VJ6�o�axK��Mb�z��	)���-؎�*�ˈRmS�"�+~�`�?t2��$;R?e#�3���|��Ay�M��~S�+s�^�.0r���p�Y��O��<�5{��	h�>
6��u�n��I������Y&��iK��<;��g���F�#�#'Z�I>�����nsD�d�����2L��W��*R��X���`z�y�ɧ�v.���p��3��[�L����ҁ����"���[�Y��UP�g��{E����������T�V*(Y���Q�pܲ�m8�2�V\P(�1mk�n�*K���m��V�}U���Q��Gv�"	��I�-�4 ���>�K˱������ �XL>֡��2!�nO�q�	Qf�@(��E6a�Vex	�d�Jd�j�uJ��y}�9�ON�L�UV{^HX�;����V�Ѳ�]�G��MTU��q��_3�L�� e& �rgm������d�4tv�]�+�	����hx�_p��v&�&����&>��Z��K��L;��m�ĉZ�J�iG�Gܢ�9
�T�}_��"����:F�;R��+FxHsbp�*_�7��EģwGwzH9������Ϯ��/*�Z�I��⾈돰����cT�ak�Y7]��vzc�gby*�7�4����C#$GqH����&/+!���ӱA!�x�{�1S�`�
�]׀Ӓ;^��bʸ7�� ���q��sĒ��Ǎ�yX�@R�F���r�y�p���~_	?�>�M��M?����[]���2�W��M)|Ԩ<U�����:C�+�8��а��ɉ������G���3#�K^~��L��3���n��3{Ǣ$��)�l7]9w2K�|�!���~g��&���\9��L��+1�Xj��T�s�.�n��=���Ωm>����@N6œ�B�n���wM��	��j� ��XK��^i^Pa�Z�M�Z�W�1A4��3��4Vy��8� ���W����ǡ#��p��w��^��=�,{��l��Y�w���_Ud�O�����[g�x�������[�����Z�
�?}�/wQ�R��с��YW�|�$�lrZ�Dnd�9g�W�.m�gws�@�9s~ϙ�z2�za�!<��)%����+���&�YG\���f��8D�zU %
m��R�]T��5
�M��ic����<g�+�pL� Y2샥$}ь��X���K&��s�_
��H��C��@�2;z�'?����uc���{J[��U�$�o	~�K8w
2�-��N��D<�����1�h�í�.�jY�wNZ2
'ùFH��F���>(2�E�5L����q�o��62��$�����~H%J��>�r+j�A���I]]��.-Y�9O�"��?�Eq��sG�l�k1yD��M������ ��áx����Ӡ��郎iȦ�u��@Í�V�kf"�����(1���5���S�$#�����cnH�F��3�p5�V�f�=�/��р����f�R,�X�����F�[B�iZlB)�S�%���U��؄����$rK��,"	4sK6	�o^�	��$��e�CG;����bJp)P
� ��V�]��='�徴�s�Y��`J�w�!�-nUku -ںS[�W(e;^����Y������o|���ɘFٽ�yG����T�X#�Ӳc��O�,:��_T�ϛ��٫�D��a	����>�7K~�V���2�r�wH,�;�^3�2�Ai:��PmE�E^<6�UP�i������܊��v�h����#x�H�:j�y�!��*3�M�)Ko�Y.���
Q�<uTE��ul��#�OZe���Āg�������Ĉ`M��add���خ���41N����^�1���\������34�hyP�GF�R�B ��56�0Z(�?8���R:ܙ�����'Œ��	�,_Kq�3Dp��M��Mm�[��Ǌ�#kL��*���;,8-/��
C�����)�(�;+%��uY:����������j������6�{H�J��{|�#WO�f���1-��`��O��cEI ��f��0k�w�X���$����52�d��L�1Π��{�	��k���vy3&���p�d�V��SD�]���	,<�){�ȶGP���W)�x���`B��km�WaX`��k�qh�������<og?gg�C)������锼W��Z��OR���>���5�������Y�g!C1g�+�)O#9���Q���,*)EA�d�,р�z��f�2 ��f@F����ãPofme�������Hf��{���2d��ò|>�R��g��, �<��S�M����p�[�iNkQfY�d�1�WpZ'6�¢��z����� ����B������4 ګ����|�Q,8��� bj�_��鏵"�O����zО�?6\]~��<1 "��'�-��_�J�zЉ���ýܧ6��M�6��mzL��)�h�Eu1�|#���KdLW"�\���*�N4a��o��P�S"�t���s��R�Chה���L��B��2��Ů�i�\�Ѡط�>{�dH�f��]r��ڙ�n�4��h������H%ZAͥ�U�,T����a�;�|�Xb֒�Jrm��>n;���J�{��;�sv�9�S��ܸ�įW`�"[ �7%l�����a��"�\�Ԃ�q|W��zif�G*�\?�	e�gK|B ��s��f��I��E(b������^Z�is�;�@^c�A�F�f���L��#���]��cW���I�GBgxM#�*�3���W+�CV�����mG`��Dz�+�,(��`c������|�6}�Ъ�C�88�%g���[K�Fɛ�T�U����m`�N\�Ј��?�ҿ/n�pR�`�愐�[��z)[X��{9�*#R�_(��<+lDk,D��>� W�fU�hY���MJy����r�oo�[��F!�ę��-�d����yq4Q��t�TN+0���G�3�k�3��`����<�DƓ4�E�o7�Ɖ�ppe��F�qq\�Ƥ��#�t+��jy*#�>W�dE�������)�-v!"�?)� �Ɔ�η�&���yx�A��=9+���=^�Ķ�1���sl��$*�s������[�8����_�U���( 
�����&W�^������Ð�r�����5p�Dv$�Y.�����R���;s��'�Tp����Vk�!WⲭR��`�t]����U�"��uOn����u�S�B A��R9H�=�=#`3�%tb(���b�aB�L�	g��s7�
��?��'G��d�zJsS����d��j�l�����4B^MئA}r|7�K��F�
�'W�^n��4Շw_�t�ù'�������{���Aq�����)d;8˜e%�*x��z����`��fͿk�`�tt���-�F%�-�︣G�����V�$�,S��t 4/n7뎉M�3A���_��;�uUy�4���Ԍ���0�O���O������+
'��V����9'	��Ϋ�%fW/w1 ����X��!7�y"�\(�ݖ˩@]e��Ŷ.�ʦջK����i�K}0e���y8���LoDr}�\�~L<���������p�@��^�wF�P83���п!�Zڠ������R�c����o;:D ��5�E?C�TVڝ�p��f��j�lt�vX���Gr�$�^2�U=�@t+C":�P�#k�#�E��_e��O93Dp2�kjO��̃=��KvS[��U�RW �Ͱ��R۽D��L�Ў�_�٪i�
��G���Ȥ4��O�U�W��rpoq)��1țUN��qXR�z��ה�W��M���J�1��q4� ���~����m�[&��ƌ����FH�ɐ����10t����UV?��kf쿠Yi�VL]ҡ�۾���OV�˾*�[$�Fuk6aJBd\�`)xqo���E��;�U1,̂�Ӎ�3�jw�d��֝`�+��Z���&ʜ��L=tG.�	"�e+�	nw�T2��r�$�aҦFX=�9i|��v)4��y���=P����]��\a�"���&�GnoRV�zvƾ��B��]*FW��B��RȵV��?��
��d���SFH�.��
�>\�ܟ����X~���2���)'���w���Q���v"J"�:�G�un��Rae�˗Id��[�I�
�����bĉ������o5�i������c���fҶ��ty��<�3�8��v�{�*v�2�s-�D�q�J�D�$��t�з�&�|1� ��n�)�� ����`6��GH�)!]�K�*8�s��4����S��t�\������(�$���0wY����l=8�9�����QS�y�8[Z��eU���{4�b(��*
FF��vŀ��=��q�V�M�?Ds�漵�`�R��
3�!Υ�^fSh��o+���ԫ:�F��gfD�H\����PW4�ELB�f�vG(��V��0԰�.m�X�nQ�N�.�D�ޜ?^�����gQ�3w����k�P��.^�n6�1Y�vV7��!��+�ۦ	L���7��|q$t��M���aP8T����p����sg���8Ƶע�����JB���><�8MW���k�6�����׺h��( �Q�f���k�3��b��E��U�`5�f�u7�k;�����e�6Q�_�˼�m=l�y;�Z�'��Vdv�<�y�<�4�����1��1`����+ݨø�U3/k�
���n�����@�x��h�V6?���y��!:��]7�.ѹ�,���3"�*�C@u�	�|�����Cm;UM��L���������dQ�����Qg���n@�;L�B�n�w(��=3<��E�jT��|������釔#L�	�ӻ�dF1�(RM[c/�v��_���䛕[t�r�<�,*(*�=X׈x4̓Iry�T�>���Uˢ~��S��(� ��*�����_zw���4�����	�"��~[t��Q=�'{>��|��tQ�4K#^��_~���*O�	-N4�t� �8m�!
����$5���@��(��1iE�7��Q�*�PlfW����1$��&'�����oJV˳޻�a��3�k�Dg�d�ᯪ���B[k�Ao�_] 8���=�:��5{D����W�h�w��7�/"p	�k�����a }��je�N['����S��N���CT�훔��>�[Z5����uV\��3�/j�����_�������є�ݰU%~�CI��bu�S��솩��#FC�ʷ�@��r,��a���
z1� J��w�X�&Ǣ+s����ZeoE��6q�v�ZR%lX��ː�jF�5k<�qYo<#Q�I�XhS��{='�����x{��o�ҩ;�Hb��3���˅*Q;���$Ѷ`p���9������̪0.�9+�O�l1:&�m:������OK�< ��1�����Zi�MiY�uX�\�*�N~�hȟb�����%�F�}_��
`"*GT.xߔ	qI�7��Ã����͢�I~h�οr so�`wp���j�*�U��K�[��@5���f�p����f�o�
7��e�Fգ=C�#���t��l�r_,zax���S�X��!���r*��h&OjDA)Q��c	�ܐ=_�>Ɇ�(�7Gn�'l3ri>k$sk��S��?�o�텕�a����IE2��q�XW<�#�J8��҈�/�F-GKaΟ� G~��W�RM�#"O��L0��>�[=�Z�� ;+�^�[@E2J�kǙiTj�;�S����$�myi�]&�j�34���ɼ-s��L��?�v��,�g�IF��s��z���;���\�*m9�J�X���%�;�رM�ݹ½;�7�b����_� ��2kw=��0�p1��Pyx6NN	�_K�d��NtMA��7�*i|�cy|���P�y�\vvP�0O�H��a!�G�%�����hQW�Ax��f6��:dͮ���nHd��#@UgC��0p�\=u#c��h�e:��!��G�p����. �ܒ����V	�[z'�*�:��}C>����OZ/�(s>�<�A�z�'_��P�y��,�Fp\���.6�|N$$lϲ�ip���ֳa-��6����������'�mn��6X+A�=)Ә���|���k��vp!#��r�/N�>��{	�3�C��;F._�v�<}k'�2�w9�l�T��"?���%��G�ݾk��!˺q>:��Z��1��8)[~5����4�qy�.z�Op(L@�5Kr��6zq���)��q�G�Z�t!ϡ��BN'Z���ٺ��	m4^��P���ԇ"i�R=b���3��^�ރ]��%��h�y�������bX%��ǁ�g�ـF���� h؏Mg\�:��@(�� �Nt�<�0WHþ��[��\q�'ڃ���B�r�ց.�ˊ��� �8弭.2J�?��k��b$��Y̓�1�{ b��һ�#Să0A��m7:C��ցy�5�>t��EM�}d���CĘ0�sNS[yo[�X�Խ�߭ep5��P�'&�������J��y�.�[�f��3��{%#��ܟ0��Dj����K�R�6�%D#���ϗz� s�����&� |!>���b�OpZ3��k�8*cp�$4��cTD(𒴤F�8�)�3�E|����w�|On���%�4���ں�*֟�}��hS�vy�Dɬ��o�xm���g��v��g�I��xW/��>`F�zuͲ*�*��"��E�{	FHS���]uI<�-�6m[�����f�7��[.��Pة�]�ZY�v$?*K��5��$��4�|KA�i��Ii� �v��~������3�@8L�kř\������G�6"f��.�u��A�#�;˷"�h�?� h�(� ��l��5V����R�]��T2���v?#�Ƣ l�����_�C�l��x����� ���>�m�CG*�A�]�����[��ѝ�]8�!����[ [92��n��Cp����n�E���ʁW�?#Qq�`;n���aÓVP}�M�<�},�.7]a9�n�h�^4q'̌~:vl\x�4G �4&��"i ���v"�i�'�<��q7#hv�ݯ�nD\�G8�P����-b�&���|�\{��/k�}�z�i��S	sA�;�mp��=���"���]T8(Y��@1����ӕ�=��{�����p+V���������7�Ϟz�AJK@���J#'�8�	���D��H=k���}�`�!^�Ii�U[���������Ci�(���+�5�I�������R�sZaM�d$�x�%MI���Y��u���E�8H�m��| 3v�ZD	�,4�42���\�� s�s7�O���8����R�9����"�@?ύ�w���� {�� _����=��a�.4�=(��![ ���@���w���GU{<.�!ў��%
[(���ǎ�`�'���c"@_R�r�d]x ��/%I0R����N׬��x���cȧx#0�]%!�����}}Q���'g�tp-�A�BНb�cF��	6� ����]�錻c�0����G������.�f���#ǟ��׭��%�%fyF�9�/�Ȓ+,U ���j�fV���WUȕk��I�U2s��h��Ȧ�ɶN?�#���8G�`�����/@��f׻l7t*M��5�2��-�'y�k�0��b�O���!����������5>5��e8�ʭ�9ݾL���"�~	�E��j��@c��(��8�HM����.�����\q#^�?ϟ����pS�����E�ĭ��*�~�a�=�#R3#��v����&^�$Ւ3�V7�Jj����x�{����rp�e���)Ķ��GP\4������(T��6	2{Q�W,� ���=�ѥm�yݠ��Z7�M}(q��[�٥����X=�֓(�aE����6��!��%��P�
�g+�f�@�]]DlJ����z�_2�q0�Z6��0�dT8P�k�~�b�H����e��}{�:5�PO�<q���2�m�D<8\�/���o���Z�����X�^�"\�{���扤+��N���M�2��ڬ��1>E�p����������C���k_����&�Hk��O�,�V�mG�*^�t�,��j��0#�Gk����:���Xi�,1V��|R}q�z�**~F��b[����P�}�#�(UU5x�C��a�M]��Oc{�����)�U��X�s6����ͪ�������өly�4Q��M(�[�F�G�q�CY�������&�).��r��h���Ȍ�O�݂F�#0w�F)Sr+A�����4y�%71+���{=��U��{����2��  L�s��ޭ�N�;�F��ɺ�D\�@�7�X���A�+����S�I"|��E���X�E�xT�����܇I��(�$�P�aOɟ�$�+=���ܾ�L�+��ٷaS6"���ʎNp��;͖/�Yh��������Y�\��G	�7����,{���|X�.�o��Sm`�hO�"5��35CdN]��x��|y)�@߻��3"�3<�W�`?a`之�]�o,0@U
\�Ñ�@-Y�0��A���A(�`����u�l�nXAr�q���o�HB��5�t$��������ǌ��8:�Ot.A����<����<�����[ߑ[���-��J�H��z4��$��i�N�G����i���'��)�[K�69A�� �k���\�Z}lw\�"w,/<�NEZ������d�g>{�8�G��r���ꩵ�����톖4�?n����i%'M>sDe�s��tn8�:�`�mrHY��(-�<�]4`��)�!P�5i��~��hT{���-0�|�����`��.d�
�l�[,Yb��[�Çp��P-eŧ���IQa�\5"�����������d�F�Xs�z%b�۲N)���;�34��2B^�]�<�i5���6���c�8��$iM�B�U��D����:��W����T
��Go������'��Қar����s�L�����(;!���~w�0�'br��J��cg�^x�LC��u������N�'�@��j�GFX��Ҽ�f�\�1kAV�>*���rI�T��df|>g�9P���e�ߐ��0Y��a�J�j��}\'Ҙ��$@#�vI��$ڝmc�V>J&
�ͬ�]'Yy��]Ӫ�?�'
��Nf�ͭg�@qq@��.m&V�[m�AP�pC*���q��b�I�?�z��/(��W�i�B�]2�4�op��k]O,OK8�&�ul��g7����j]HJ9���:Թ�]��:v(��S�-��T;����;��6������ 5h>�Y�d�;�7�I{�	���v��$2�
ɻ���~��]�����!B@f�\�_�E%�j<=xsjO;�_0�c�)�__6�7O��>5���nY����:�	̔-?�6�IL�G|R>mp9�ӉZ�(mk���چ�C�>���P����m-g3��N��Z�Z��o�����:E�t��=��Q�+���A4�z2���'�*B�Z�j��	�o��j�z@ǥ:9[��t*���*@VQg[��1A����'i��s
Q	V�`c(�QFN$�gP�F4CI�C���&��y�p�>�\^t�sۄ���3���j�����F�՟?ɖJyĸGNߟQ����C�[A^��Hxvz{���Uek^q��1�5��$H �
O����;C����p��у�Ly{>��K���P8�J�=�Sի�ב4-��[h�4 ĭ�Ka�u#��g�D \��@L�MlƔI̣������c����f8y�K@v�>��ѱ��ލ�d����	�mQu�c�u[+��&�w��>��d�h�� >�|�v��e-R�(;�|#��-��b�H&A��r��M��{DHzN0h�E��~����{#�UA"�ֱ<+�_5��j)��[f�UF���kUVv���,O��a�Mp�a����C@��w���<���ԋ��y�����|ר�G��xI���on-���M������cﰪ|��f�皌��3t�{pM/���n�($%��?7�h�utKpY�d0����(�:]v�Ԍ�w��M���i����7�����b���HԴ�UG�Bhm�f����Y(r|����Y���������4\�
�1��\STQ�r�A&
j���AC1�a�Ö���%>U���&�0"��-, ��-�5ӣp$􍒮��:�� *�ja�*�O^��v�4��#�R�;��+��Ҝ.bd*��d;L����Uom��j�"��[FӒ�t}KI:6M�����3mr�\7g�]<$�C6hX_�S��8ga�VT�'�V!+�M��y��ЎQ����Č/��N��>�e�N�gOF�i�V������2�K���`ư �#��ܤ�	�+/�Az�ǖ��.HǷj�yeM/'z�'8������ �y���4<��\��g��N��\�,�>���-u�&�@���ЀƝ/`G���?�~wv�4���A
RI�z	�9��,�E����K�H�5���PtkǹU:�Y����D��p�z'�s^��̆�/�_]���=�ui*�	O<Z�Xz!2IA��ߥa>n꺋��i��u���Y���c4?��� �י��D����&.Wj�!��&����șd�K��ӯ����!s�S0�%B���Z)@ѪP�!%�T�F�9O���ԁ��gu�~`Q�(�b��h�t�!0�u��
��	����"�Ǳ�H&����Q_	R,��*���O0K���d�Y�~N���7�ݕ"Q��\����i�ȡ�������ջp��#O-�%����6r�WX_&���7+"��'D�{���n�+/A��B�ՌQ������ .��3S�̺O7 _�eȅ_�6���m����fok�.0���9	:}㥱�Bs*�,���f&�t�9\ܶ}�a�K6s�>�'����xb�ZQEc�'���Y@��L��%��~�s^7�2�dA����1�h.�s�]��+�(�5��BK���I��!��C�t���I)�c�0�ݩ�B\Ĭi�t��ϱ�MO����C��4?n/|��~�y��Dn� �<�RaX�3%q������@����t �W�1�#mX[<�{���^�␯��#��[��O�ag�]�d],�0���!K��)�8EjN.����@nǖ�n�([ahv�Gdj4�3�OS�>G1D���B2i=���!p)#�*�^�̎t�
C�ާtD�2�#T��"���C̘�н"G�U�*�$�K%0���v1\n7T(-=o�W��i���LY����f�o<r~w������ee4��~����d�ZQ���^C_�.3�W?@�h>D�#�V�p|�"`q?�'�^��h�%7/-�f&�� h�^h�֬XM��K���c3����`W�zxm�U�Dy췍hb���Yw�:�;�z4�I97NI�f�	n)�ԍ3�WRE:��c��`�V��=yɀk�6�[h�Ѩ��z�ۧ�B�"& �8��6�4=�WJّ;�&���1Ċo"�d@2J�p�T�uK`�G���;O��]}���[�	i~�Y��e�����oꕗt����!��j4(P�+3�Kd$њ��z+�k#�h`�.[��� ���(4\��a�iE��6y�+�N�044���ʖU��û�n�������2b��C_(����S��!ꁡj�@�S�~dD�NF�l̝Q�h�� ̔Ax�C��T��'%ؽ1N�2rPP
���}�$��s�Vt�LX2Yw���vC�즒���j�5��M�#�̔]��ieGw�p�����`�7N��t��BgS����(aR�g��Np7�I�n[�d�}��rxò�l��1����B�,��
��H��w��o7(7R~�
�ٝ��»����Z,���U�L3��2��]�L���U����2�͇��؂���[��R[�D_��q���5��(���qM��b�J�{�"�/����z+NL�*��Y��ª�S�G�Ĝ�+9g����z��sBi��Ċ��8�-��ڢrLA{��jviK��kea�s�*�⷟��c�Vb�b6U�������a8�Ax�x��c2�b���s���렖�I�~��0��/�s(��r�i^6J\�י�U�wt96V�g�=F���&9d���[�O�ר�;���>K�W���4ʻy=r��Hf��ɩ��Q�	���dH
��fV�_��sD����� С���f������"D�F��	��ʈ`,�Z�����u6���E)�v�EY�;�	�?0	���䪏���m�~m䧉0����Y�-p���'��;50
�LU�#���5��'B�w��_x�Ho�wzb�>i/9��"G�K����/���oE�d�@�	_�A�¸k���i}!'��E�K��nz�8��]�h	 ��z=q�����>���{"`�'2�>?�S���qC��,v˘�����6�����C��)�o�n8��:sP����e��#�D��y$�|�χ��D�*��N��?���!�\6�Swa���Τ�������KE�4oϘH�f���'�̰r�3}�N+��R�	���)�緙���p�Hq���{*��*ی�Q-V�u�˼$ߩ_�q>&��9mlݡMݴa�����kxI��"Zzt5[�3M�����i���D�Z��M�_#/������oy��)ڨU�@�Pxnᯀ$��A�T���"��y���^�#���OKb�2���
Mk��W�AS���u�y�p$��Z2�_��֌oW�N{V�=-�&-f �vcì�f3g>�Z�䞹��A�g^]�-�#a>�K��\��A���p�d��A6�bq����pCB[�MTXr�4���=�Pn6�S��htT�?==�;坭\H�7&9�����=Xȡ�ʣ���ţ�ϋQ}}�aD:�R��4}��i���v ;�,�KάC
:�|�د���5Er����U���1ʝE|��2Z�p��W�zG��g>x�<fa�u�{^����r�*����\�j�y��3�U/цrg�R��HB3��P6MK,�?>7}���23�Ȇ��\o]I���J2���f��`��ˋ��!ɑ£_-M���]8Ar?���%J� ����u���5��wz[Bx_�03Au�ϸ�8�i:��V��4�6����Jt
�hc?�9to���c|JFS�LU��T�`8��i�@����Mv�Y-d]���U(�]�6G��d,���R��'�ҳ���P��U��o�9���U���E���zG�<}����𾫒q������G�oͩ��0�͠�A 5C�\�PGqW-��}>X=PiU�@��p���P��-s�mt;�PIWT�3{��1��	
�LW;4��%����3b��_��LY�.}��۱�j���s�5�nU�c[���@�n��c^|>���ej-��Y;�z	�ƴ�{=���Ҏ��
�x}�ؾ���ʨ4ޙ_���3������ ���)V������^^��ϧ����$W
|��n��}���������=u�b Y"I=\{�H�\_ ���9&���\Uy�ZI2?����"8�­jO�7:L���=k $���n���D����:�O����:�iD���N-���{'��A{)���:��3�\FV�Z_bRW��1����y �q��2�p��$�U�A�m�q�y�
Ӣ���p�c9�:�xE��F�V����(��q�H�o�����(�s�ԓb��e��RL@�� �T�p����߸�o�E:U���*�- ��,v�h?
÷��+q��2ˉ���!��ƺ�=r��q��Z����bAO)��'�b:�{.��<���|����k�@�r��"g��C���ZziE�?�p�)T_Bl�ԏ>�  t�z��0�D��ÍM8�>	w�L6�vy1�-Ϳ�cO{n�>�ڧ㳜�I.���)�R;�'�����H�����߉���3ԍ���̐��#����S�m�c٢�?�ss�f.�=?(x�;�J�PM�3���@��-��䎚��	Y��y@�Ƹ�$�)>���
C�w��(kL��|ewov�w�l��D�7}�>s
'.���36{�"��g%5D�HN;l:Զ8�cԐ��͡x�B��Dv�s�R]r�ջa��F��~����C ι��Nqv�v��o�r�%���<x���'�4p�T�?j�c	��h3�.�
���9y�"MHp�X�H��EY��Y�&����,���kq����5��7�Kg)?� /���E6.�֙���w_�2GX�S�`��]�42��B��i#;�B�/��i7���Qzzġ~�
�ѣ�ϻ*��8�������<�S��$�]����2�7��1�'<�L��U
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n�sC���}�z�%�������๰#�1\k�3��p�l.msxוYv�m�0�� �[�T4x�K\����M�\<�q�=�F�ѮQH�0iNLsu�P�%�J�^֢�k $��}�����d����M�k00N���)��8MM��o�'!�r�
�0��"
vW'4���y�yK>yl���o���������J��Ϋ�����dW�	�_#w���������[=׍�XT�ȡ�rhX�����(@��e�2�B7뽕�r��<Ƭ)]��W�|?�D�B6�p����C���\���-_|J���b�6j#3�U5�n��=���.E��A&赮޷ �5�=La��A�ՖB�6����R,o*��� m�ɨ�|Ų������ֺ�g��y���o4S�5s��FaoHj�/+��!���h��6өC"��Z�氉3������('��1t)����dVh�O�������Ů�6���_�v�R/9m�8B*��c�L:�9�d��x�A���"���j{s%�sN�.6>��;W ��7��y���L=�M�Lc��*��q��{fd��`-�	�S�Sͭx�p��Y�,���;+X��[<=n�ޯ��)[\VV�}3Ő��~�=�jk�ԚLh��Jg�0\��O�nD�z'%i�������$@+�V8���������{a���-F�Nn|�h҂�/�Zc�1`�D�������pIy8VgS��)B�J�K*L|�7�'��r���R�!;5�xI?�J��FEr��E�#Ux�9|b���D+ov��A�X�f@K���uo�x+�Ȃܦ�.��?�Gq�a�aN��S)2�Z��Z��z_��K�Oן��!&�X��Ff�����s��u)Q	r�����*]�fd�q�����=|�7���`2��Q�X!Y��K���J띶��Af�O�@���d�^�h�I����1c>UWy��í/��4I����� ����`�����`��۲��8����p^���$�Rv�62�. }`@Pײ�� 	�B�Q�,ϰJ
��\�&4�i�-BߗG<�P�"�\0�����5_�	
�E+1z�|���1s�K�(���7k�F����.�%U�Փ3�q� ���h�Mb��Mq��Jv���9�k˄�_�,�Ov.&���X%O�î/M��{��h=҂2�0H�����C^h
�[1Ǧ���J�i�vy-��k̮�_��E�w��>� F��G;��oa�$z�-%�b���i�K����Z�:[e^Ħ�#������J�O\��(`u	����>p�/�7Y�Jݜ�@�?jkAl	�qdb)4���,��}�9N��'�H�.��n�����XՅ���#�׊66:�_��m�V�9
�⏊��G:�Tp�W�C��Y��%Yg�o�� iq,�/�`y7��[�۸�H�-��'X��w(�~�3�PҟE镳��P+(�A�!�U�4�|&5p(����oM(�[���)@�P��q!8��L��d����|ݫ{�5�36��)���#��/��r���Y�J���y�A3���xY;
�F�)2�����}.	�eq=������ ����xԚ�5~����|i&��.�q'v��'�0�k�{d���462�j����ʅI�Wc��eR��\cT/wb��"?�Xj��t���z"T���
�G��P����M�k_x�T�X���%���?��-ocys�b7�^��s�Y )��/��$��>#��#Q� �tg�Q���얦N{}�{ll6�!�]2y��nt��3�6r�ga���-~CK��P�1�űXNT������S��/�;	�"�b0Ay��	��%]˵��ŷ�F7�\���K�����_K�H�1�1�AE)8�$�ǡħ $�G!�DiN�)=?�>���oM����1W�&�T���J�A��2�ҭ�G'%������Z��	t���0J�)�o`lP���o�f�z��k1%g��fp�#����WéP��2��Z�`���k�h�?W,}���Ͳ�O����^X�2�KJN�uT���Eo��ą�qVL���wo]?F��|)�
h9x��2�&o�y�C��caC7��w��U�ޣp�g���~�'�fl��N���:]���ɨ`J�)�c�IT2�aԄ��MB.�(�SĮ(�	�� |�~�	�������d�ϬN.qTf�����k�e��ݹ�=��~��;-�k
�[��5�q��댷q��K�m>����Ѕ�v�T1�(e��K���]�$q�?!�@�BE�8eaK�h����Ub�����w�H�'�D�T]��q��2�yw����`u��t�@�fB��S���6M����Qm���ނ�:S㩊���Y�������J�n��_�̓2�(����0�[�B�`�p^gᱹ D�R0��!̑R+��:�F�f���_k�R���T�fn�c��Տ����M��i����=���t,e3�"*�w/8%�D�x����[F��9�M�oQ|Svݭ\�χ��*�Nj���c)ܶ��<����Ag)$}�%�����iǚQ���p���hVH��2��>��o�A7p�l-��׫e���sEM��[�M܂_�ײ��r��(X~�ch'������7N�;qv? Mѥt�%h���9S��HΒ{w�������v��D�d{:|Tu���:*����ˌ�Cyz�n�[��UzS6催���	�{i���=�P�(����V�����{f��bk���>|��}~�X		�-p�9��#�=����Sf����&h����U�_�n�@��7D]�}�N���Ԙc;F����QkK�~��,�`��c�H �!�7��6�50��LQ��@։e#�G�~����?�} jSG"r�*�o�/�+��Veg��،]`�GaK��l�JN��	���]�U���a��+������=)��i|��[1�\�:�rl{l�M�?�0��:[����Rw��Q��c�a���
�Sj�ĭ�hk�0�׀�#��KdhH������~������cb}��e��0;/1�}ޡX��[$�%��CH��Y��K}�V�<l0A��AY������6V3q;�g��~yq)ô!�\7��\Ӭe�J�Ȃ0�;- w�5�%s���[��7�Wˡ�R��_��^l�=��;��U�Ql�B�6����P[�a��tr��/>��_��Kď�Y���du=f��MP�T����n��"��ѯ�5&���9��B����Ι����R�o����&}є�+{d�a��Ѣ�?��2{���4rΚ�s��� űQE���c��]��l%�xw�u-���7Ps5h /Ղ� d��O���v��U�̌VD��E��d��4	D�&K6��WJ�[r�Z4�E�n�O�I�SP-������ޑ��̠b��*��:������H!&M�9�����Y,c��%WY<]�54��8<�#7���4+��4"u摙�XD8��-kb�V��9���ЉZ Hð�ĳ@^��H�v&%z���'���k`�}JiAj+�M]���J�-T6rq��A�6�t#��a>u��(X�K)�P����$Bę�����y�³h�R䝚-�J���~@�oB�a��Ca�����f;�����F�NC���oc!{�|�mI2W�s`���0�J�W^�ř��v���/�{cݹ=U����� r�wˊЈkb��^I�6�B$��:���Y7p]ȕ]�k���;�}Ovh��P�oH����� i��zĤ�{;�|M%:�����`D�\3~D�0�TTs��:m�3��y~Pk�B��a"��#m>�܈ʯ��&#cd}�8����	��}9�ũ]8r�+YV*���׺��
�2�����9�$rU!�vM�=�(���=M�e*$��j�A�E� +E\�3�f����>w�[a!#I�a���!d�8����.�o�ߋ�zӒ7w=�����x�E�ۖ�k�+�x��{r׊�(�2�v��<*�b�6�a��&w��F;�*/)����KVF���fr<Y�e�+����'�I�:� ���8�.�Γ���t�K��f(�����QR�x�n��[z�������{��[1�w�]��a�>�﨧By�b151{�+P�����H��_^�l-�Rm�������@�u�VR�9}�(���<|5��X+J��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf��((�yH������Xd��X��&M���,�Y�h�;�:�ɏg�a���(�F�� 6A|;Ӗ��'���nBq�r&G7�ל4��6��1�]���u}�Qf3��/���5�-ބm�7h����I�r��i�*S��Y^h
���(fʱ>I�y�g�rso�cW�o�/$�A[k;د��c�b��M���E����g��� ��DkgBU5RY�6�1�)	��(T�����r{io�%�ʹ,`=e��C �3{��U�Vs����S�;]D4B[5�v�Y7����:t���Mz� 	$V��~�O}F�CD*�R�~\�3�����I���T���{M�� �ԙ���W��\����.������&S$�ណ���$� A��������R7�@
UW1a�������Ӣi;=�JBL�怤��*(L�^��] A�����[� �m�e�f$��1�|x���{@���f�A�*ϼo�P �y� h;?��t��pk�_8v�����D�������r9�9;q��sp�������6��Il��"{0����B��$�	����w���c����B�(Ԙ�Vq1D�v����=��<Hu<zH��.�^���.��le�2�<�+��{��Z�8Q/ �5�=%��;.4^��x�U�jNK��VCP�����K~����-�4�R�~���÷x\~�G.P8��%�s��~�.Z���5n#Uh�P��^�r �4uP�<}�{��]��x�NZ3gD@K~k�6�=�?[��83�򗧉�-R=i;���Z'Ҍ1�pU�q8�q%��w+e}�*��ў��#(�%�@��K 3��V��6�HБ/���՚��MC@�s��+�h���T�U��)?�.�<���Jukz��6fo�kR���CH[�p��g&۪�y�˒��Ɏ��^��H:�t���r���ČP�U�35\%5 s�ڞ��Ϟ=e�V�g�-��u�)�#^�5�m�d��7�{�N2�<�,�/6|{�ЯF����X�x���	~�ԾI���;G���[�l�ziVtI�b�g~Ȳ�ye�t "���$��)D�lciF3���{��Qt�;+��p��b�|���|@�WC��wsq{Q_N�@����κ���i�DY��6��r��tpO�M�)��Z�('Ѩ�_��;�O����ҽ��[UC�����k�}���hH<= �E�!�W���A���Ih�[���̅4"dFmY���M{5�������|����Z�t�G��*��1���4�A7x��1�^�c�1c2��P�v�Ҡ%��iF��Z
K���+���g"��eIv18^�h//��t5�3�#?	���eS�o}��	Oo=�@YU�L�[:f��jH���x��,�td�ke�͂sA��|��D�U7�\_ܲ���G]z�ߙ����k�	���q(�*��� d�aR2%S[�t������å���{;�j&�7<Xf|�o���d{�u����ݱ�W��9˶�s#���d��5_�>��ºF_�:�Ŝ�[Xb;�ET���,`{�f	`9�?ݟI��b��m��; ��s��&ڦ<ō\$zx�f%_�5k{~�NH���<
�ʊ���,�*�]gf^�=A��&�jPve�<;��f��W��3��GL��L�g��c
ot����L.�(�˵a�9���_W[�+沄�G�^��~3.-|��a<� ���|�k��Z��������;�,�H����Lڤ�y�Ve�����I�r�[S�L�7�?��B�?M�!�w�u�_.�#���d�'Jt/�ׯ&���:�2(3�ʶN4Ġ�J�pI�޵�_��ks���ыi�FG
:\��R��Ȁ�g�o��꙾I��(u^��Y���ա�j�ɟ �V�$��
��h��({�0>	�}�DP4��L`a!١�ƹ����D��U �_�9"�.��1✢yuÊ���������GN�uA`T"�5u=�}�G�����w�
3r�>�IW��̨�k�k�
~�h�DH�&��!���a��z��mU7�����盻L`9���b�B���M&貳j#@�f(�M({����u�I}���n)z�ۮgj�G�t)�3b����+y�I#葉�x`�r�ǝ�Q��M�y��4��w�_D���!)!ளpaa铐�	E&�G�#��(�h����^�g�Li��^P߉838V���*���r@��X�Y�|�i�)�L��m���`{���A�J,�p��5�A�ak�� \%���<��)DG��Y��
b�jKva4�ܦB�}�C�$��5����%G�gWN/��Vsi2S�[�ć.� HN�&i/H�C�49�X��.a�Ȉ��O��l(�߽�~�\=��%஛�g��t���uVѓ�'�n�U�kF�Ɂ���H
a M��Ub��னEF�i�~�X���?Z	v�ؠӓ`��Ň���$�6Ɩr���D�?Z���3y��<Ϙ!FC2������9`D�a��D�9oؿ�7����.P�0�n�"Q��K�3��[��1�&PT��)T�	׏�X�}q�q%��;�� Ó�.���Ů>�[�$���^5�E��JΦ�����j�m��/r��g$��z��}z	��򰽝�#����m��\�ʪ���Lc�E��¿$�����@���(^�ְ�`�5R����&�  ���l�m[X^��_\xȊ�L�51FGq=�,�Jr>X��D� sI��ۛ&�<��C����2��c�c5=�3� ^e$f����N����b�;��A��,j��Х���쿉��^���q�ہ��@�(�=�C��vE2�5tw'�⭍���⁋}	߀���mm�bN���\=ϯUC��zZ��P\�8�j���3]��<���Æ1/�|�,'��T���6W*�zdA��E���N(#��9�y#.��_/'�C����^zAe%�z-<�<�#���ǃ�ص�~��L�ܭ�DlqMӝ[��)�4A`*���O�=�����v}���G�j�s�L�;67���)��b0	f��g_X�>�ϪG9�"r����E�YТ�{�V��{j�'R}����$���:#�Ȑc$����&�L�az�/���7����a��\��8�C(�A;5�I�gC�`�����3K��V0��R�7$�iӨ.��̃y���D@{U�%���>�`�G�tH�{(9eP�_2��R
��
&�н�̏i���&Q�.�c5I[,�39}\�q�	��y�����#x�pl!�}	�W3�Ge��30M+g[��W�"9�<�J�~fJ[���BI�*Ė��VO1޲���>�o2��GQ���]��oE�[�	UcfM�+�>Ϊ�R�+�C�e��ϒ���\f4+�!CY^<,�<� ��ۣ�Fr��<}6������@�:��Fg��}��$��]m�[9�S�%��\���W��?���UsD����Y>�w5}�_�ގ7���U���=|(����?����ߺ|�#H�F��5iG�h&�����3�j$5�2���R9D�KYBw� ��I`������,�/��3�6�Ǒ�x�U6�@��9��b��7����d֓]AZR�Hf�;�A��n���$f�I��(^�c����K�!�z��&ި�����p�Dw��7�!XH�ta:2J��n���}a�M�l�\t{�����h8d|0.�&1��[�}1q�qa��ɷ�OH�g)�a�R��P�i}���"=�ǍĬ��&��,���)M����r�J�8C��
}�T�N�G��o�f�ox;�}�!��2!�{7�W����bRIs��bU��'�>*��}�Db@s���5�$�d��Wݶ��]�5�V�u���[�n�l�d�f����2jr���[��b���U�2���R�$����4x��W�AI�|���H���3#���κ�Xؘ��9띘���z|��%.#��$ �8S��s]l���?'t��S��<8n��tN�J�*!}d�����@��?V�a�4
S����u�+q�d���&��Z�j�B̀�9�*�Whq�����xY��׼��dD���w��+���Ku���9�@���N�Ϝ󠷊��O
rN��Ǻ.����-2�jB��R7��&�%�/
?K��q0=�RcAP҈�Vb�w*S���+�pv���/���Nϸ(�J��L2m�ן]���O}�}~[�]]�#Ӫ�4�F��]��lP�]�o�]�U�/؋�-���:��Ś��#��I�/��|�c>p&��C�����(�1>g�%w�����?|f�D���ƪ��+��pǰ(bt���N��^Lt��'��'c�� ���Ej0�$��J�����y~�S��OP�x>��]�.x�z���$������� Bw�/˛-�L�M�$��eR۵/��უ�*>E�N�{�^o(	���=�@"�5���10�ys�ęd�m��)�W�Wm���f`y��x���2�hٶ�^=��ׅ��,�w��A���j�PEj�I3�Ot찟Dm����&�"4Ɵ�k3��"|zv����s׭�����wr^9���8��{Ry �x	������a�����h��j��Z��3�9$ε�9N�7Wɦ5Ѫ����r0S��L�����0���g��ka��=l���Ԕ��0�$(�<�b����d� �g�l:56�����&/��.]#^�s[�$D��a7Z8�8�$�7G۩��ʢ�ħf���yrQ}`7�B�`A����m樐m5���2�%��>M�i�6�W��7�`g�`7��f��/�v�"
7����T&�o���5~�C�`�Y$�>��=��f�G����rԐs��}h$�pdI��9���� O���Z�i7\�����IS5��,���o��������p���y�.O6 ~[��[D�_��3(~d�E6:�$�QV�cW�%I�g����F��v��K�tS`\�9gW�(m	�S_pso�8��wE���4#�cBh���vG�2��������4�*�[���N��Sx��5>8~�1ȿq���1ap;瞁�{��E�F� �<wq�Ѝ(�b�i-�엝�s6��IZ�=�
9��Ri���,#<u%��Q�l������3^�dI��6RM:D�B<s��.06Y+'��R��s�Đd��O:���L��ԕH�
;r�f�[�,�Z༨�kn_lj!/B��zw�h���E�"2U�%�Z����pu�~����d����e����	�eȺ�^Pq%���J���&���H,�9��*+��d`x�|� ��$��z=�9������Qκ�W��xv�kaJ=#y��ZZ[YD�:i�,s��~)^�Wě���H��^��pb��ph���f���v�^���� ��K�t��)OD#j�SŀO��Z�ѥ�<�)f|+���C��!�w�7�?O"�������6j=��!�<��s'QGeB�!�} ��������F��-	F9�:�����V���2e4y�O��8�HڪT �вo�p[<3.�Za���	8\����=��RBTr̙&m�qo���:"Cyr=�!%s{�B�����o:\� R��wRײ/l���x*�.p�k%����E�"�o�\��O��D?�]K{�`a3V�μ.�i��M
�`��c���@.��@>�p<��b��s�>j�u�ee��Њ[tʯ�T�TH�^I/��4R�.���>�S3Ś���b�M7r��㼜LN
�Bj�(�L�G�խ�ig�T=��#O�d[�s��vNr���`���x+����I�Z�e2���
p����P)Ō��%�?�kS����k'���F�@4�:)�( ��o�������S�݆�yw���a�M�~og���mI��I�l/���:��������{ bԺ���,�ab�*�.E;mF��t�Eqx��W"�����%��j��[6Z��TG����C�h��j�t�H=�������=�T�<
x�ni�_J�]��cZ��R�B������h���P/�(��qY�_�6ۡ&�:u������ʀ��g��L�O%��Q�G�ؗ"m�SFty�����uV�n-��,��������JNGU�먼���uu�жrǛ����=����V�_)Z��,`xcJ{��L�CA�iI*=z���B�YvPt+�`ז	U���2���1ɞ(��=�L�v�~G&�
Gu�,��5G�\����Fu��2������=�^����30W��m�J��//�Jc��P�\+u���Ed�� �i�Qx�H���)1���2J�v�eN�)treGyߗxQi�M2Ջ����[��R�ݥ�{���E����j1�
 �@xt[\!|�O[m�>�o�z.O��X5��0����._hN������Gˁ��ā��L\�X�(���Fe�ٳ7�����<���u���BHa������ZĽ��w6N|t��h��Xhr�r)�m�Tz@�x��o�#gl�B�*�����d:<h�;��@�С_�2,���ԓ��,��L�֤]BUmz�N��rN�|���&����6��M��-g2l�b�S��p���E��$/��{�F��t�x0�:�Zy�.��t:a2"�u<6��*��q���!t��[l�����>c�����ܹ�j����\)c�a�A��om{˶�>SZr5�(�ғ���
@�G��k%��$b\ `F[2� 	J���Q��	U��>Pf�솛��!�6Җ�qPU��Õ��0�x�r����/�,�u���=����c���&��`�wlrs�EV���N"1��PF� ����i���g{
��?�<A*T�Y���d/A����S�x"�Rxw����eo<7�Mڲ�Z��h����p?�ʴ��+��/�9l��v��b?�
P����d�_,,�:*6U�u�p�D���a|<	����%
}�Qy��*�JA6����~ৎ�oP��]@K�9 ���xR/���?�w�-[q.sp��@ۘ=�#?L�{�W`�O�è�~r!PoG1�����
KG��
���,�r�+b[�kϜ��*��vg�⇙E�n��B�I�N _�<u�T��L���V�
~����g쓞{��j��:�lkh��3�(������o���{
В���V�ʯE��E�@��Z�L9��ZK*��� Bq�+�8���@ߕ����&|upJ�����>��!Zz��R���(����&[���P��(�;�W�C��vWaݤ)pj
b���\�����U�@6a��i�cjs�`��0��d^����4�iL�.{��^i/P�����뾄V�cL���]�s. �����)��)��ǻ_�o�ӧ];�dT�B��{�=|·�/�+UX�[n�o��X����KJ	���C�]��^��� N�%���K�)��u=�><�kb ��v��vleod����a`�b�iY\�&^v�5�ш�:�&rLq݋6T�I��xc������$@F��C}LC�ѧx7H�E���~M����VbZj۞C����>���3�͉s�k'�	a���%�)�7c�L(FT<;��(��53ˋr���J�h��T	.u��W�7��M��J!Vn7zO�&ޑ��g�!�#L���/ʃIG=�Y�w�N��m.y�%!�d;� ə��ri=\w{��s����O��~T0�)�5�r�v(�&���^�����?p��[+��AD!�a�-��C����4$��96�"
�bu~�%�^e�F��%O��+�V��Ůr���iyM �%ӳ������6\X]�S�4�b�˫����)�+ 	�ݧ��V���yޅ^;����09Z���6�{��F����;����ju�CeЪ�!��B�n#=�|��'��dd+lb���5%�xmzy�4�1]	+%�f�${�y���	����,�6��Ɓ+�T��H�n�W��׃֮�K���u�X�n�um��Y���9/:�_�:9
&w�tfԊ=��v��,)t�(u�E��.X+ʫZ�����T�Ju���N6׬u�_���/cv�¬� G�XJ���CL0�D����^3Т�Qw��h)�� ו���;%섓�7B����
��<5�K#5�YB��y�no9�@�Xl�x���YF(3���/��(�g�����4s@��W��Rꌱa������ɐ�cB[�\ 
�W.�/ne�����dF�O7��3�����X�z����@ t�:*��r����
e�;i된
>%UirS+��~��Z����M�t�+`��Y@4�/<yi}�a^*99���N�s����Hɡ���(�a �p;�uq��[��p_<��E<D]�=ţ�5�D�"U��qBQ����a1y�&��Ϡ�VZ-�G^\b6�+���1�К>��?؍'y��-S�� �a%�$�����Q3��� ��2��Bq��3^G�����>���ww)* �uث&�p�0V� ����*���\�i&�j��^�Ɩ�B�Ɵ �AL\N��ڇ���")˰ ¯N�yB+|&X�_ӎ_��H�`XYH>7q�$#��3�6'�z!$i��KHM+ӫ'ѵ��7lR����F�(^3M	�[�7��J��	�Q� 6��٢*�>mWx�d�Ӳᆩ��P9P���`T��#�>Z��d�n~s]�A׮���X�
�� ���Fr��ɉ=���2@���Kr_�&&08ɋ�7�e�����x�b���<y�T�f[�Eh�[<,/�RL�5��������ɾ�EL*� &�m����6	B�|3r�gǮ��5��W캎~�j��5P�����k_:9�h���K�A����0���p�QV���J�x�e��h�dVI2]�����q����c�9�Ѽ%�����h�����sh�+L�������q�ތ��v>�{��+}F�0Q��rf�ǁ�K2�G&��)����|[~r�Ga@=q	�԰���-.�;�q�F%Q�H�ȋ�/��<�f����,fR�0I�v�ɒ��0�n"/4� �Z�Z�t~E�F�m�ۉ8.v�z�>��P!�꣙"�6`�1u�
��J������-Rtjާ]/"�A�ЫhMm��^=���ˌ�J�f��"S����!�d��U� `|�A��q�,���k��]K�p�%B��W�3���:��s�Bv�Hc���0kMA�"JR��w�l�ĵJP� �A<ŏf~c����O���Ь[�I+��D�(`��L6�����Wb�{�rT����򽼪e�Ì ���%s�im�ưR�V�R��	�b^����}��'��/� k�L�ceg���b1���-+Tx<����R���"H�xŃ�2��bꭑ�^�v!��������h���:�B!��P�=)}��i�P�V�m�}���{ sd���MA�FNr��y�;չ�0m@���U���mW��H�/`�D�g��F\����z����%������n;������GO�+�g��b���iI�������9z�hW���!{����-�VҶ����u!rf��}�ɿS҃D:&�l���A+�Ԛ��|�������eM�R�&G�g�ԗ�5鲿վ#a�6�п�@�%�H�������9�x#Dq�U�Й��~l�8`��/T������bA���6
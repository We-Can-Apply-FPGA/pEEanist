��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
���[p�Ky�-	J�@T�h��g"���Z�YC�X�2FS��Q{D�H|���ʳ+�9�&�\v�C������7ֈ�c��/
[9����@&q8|�˺2�g��`��\�v���j�@ҊX1����.�"ci����<,�J�[����u��'�8�Py�=Yޗz�4� }� �� L��	��&���|����)e�,6���<5Pɂ[��|I.��_[��~	L�FgEBB�롄4{�~й�E�L���_,�m}�i4�~�9|�
q@%5�փ,��ʍ� ��:���[ޏ/T9��X&7BR� �Lj�����u�#�Ӈ��A��9����p	�J�o��7�E@���/GI*6aF�]�H���ԗ��J �6ńV���ۉ?��9XL{�I�u�d�>Q΄w����.|�.��_f��Cٳi�k$HZ�7|ߍ����Wf{̻�*Xd��O�xY�d��z��\�a�N�&�終b�(!�W�:�4DrTNMR}�'��4f�6,�BԳ
)l8�40�6�&��ng ���h��VQuZ!}3ؒ�~	�X���Y$���H9�����ujӓ�]���/d���ͦ�S����H,��P}6�3�t��\,>�Ҡm�O�W�)�)bB��tS�ʏWk�S�h�����b�� V�"��^@��\��ԁM
C��|Xu/�=�O٘�m<#F�"���1ӝ���4!�˂RK�Y�O��I�n�6h`Slb\wp��d�-��,��J�k_[MH=�s;G6�E�k�Ƹ�<?��%�go���)�S]�ΛYC�$r�6�P��^E��|�<!�ֽ���@z��-U�V�(�r�i�L��IvĂ��}��j��c�T};��:Y�ɊgȔ���_d	��0�R���Y8I{��^��%t�ӹtS?�3��}�_�����~�(M�r]�����~�rP�R.�I!J+�͹�M�7A̵�=hb䟪3�<�oBq��׿�gy<+�U�L��Q!p����Y����}��p;�9ܠ�z�&$Wi1��E��B,�	J����Z0�	���d�)h'g�ί����17Z�O=�O�D�J��Np�_�
Њ��F�s���I�Λ��O���������T�l(�c��"��U��f���q*Ɏ��kXy�����s�&����=L�� �Z��g����d^Г1��+��.���i��&�����5��;� N�;�3��%�@G���%�5��1zhYι�ݺE��t!�Re�A5�<7+�T��G��y�� �5�	6�a~n���(;kVq�r8��9H?��_�$�+����*���1���:�F 9����ǖFw�M>ʬ����=�POU��D�-�[ �JF��OC�UőE������9H�H�������2���?����)G?�߁^��N���� l���8�}�y3��\�Ө���k\����nXR�0i�8m@7�j��B��n9�XT�_A����z"W>��	����lsLn���*Ү��萑Ţ��WTO�r�-��;�DQ���ld��b
�z�7�Z6!ڟ$֑p�`��Y���E�x���@�H�~N��H���u�����k���Y��8q��{�j���r��}�%K[(D��C���(��k�!���Bhﾆ�VME�W�c�����+xg�Q�t��.��bjʲIF	�v�����5��&�CCR����?o۵26� ������@?Kr	HK�F��i"(JQ�EZ�v����ы���T��/���!d��AI��o.�/x	K`�n�4��2`2� �a)Ձ�#g@�5O /���?���Q�/�S��D������m�*�
���R��
v$��͊9W"�5��-�U^��-�D�"ƋbU�Ý��L����l`� 8$*Y��Y��\]���<�^#�U�v*��I$���S�DV�z�2U�-�<r�r���Ƚ��U�t㻼P�ӑ�ن��$ٱGH'�����\��)԰��@�{�|���P�y�Kc�=ìP�L��)����w���+��84X\�dI��Z��7�#:��2�a|HͿ>S5�b1�����EM��Ѭ��� ���kaQ��\�tWDdrZΣ�I��\���;ϣn��QeD׺qs��-֙�p�"�.v�Ã��i����G��K��D��Н�C"�:�J�B�+K[L�8�9?��":�a�:!a�#�dT�A400�!i��I$)]��+��]̩˩�����p�)�"��j�$w����;�� �`��D~3��U����Z�%2]M�{�"�W����-O����ԩd4$�Z\P�/�y���сs�V�K�x�4�?�9�>�d� �qj���'x��b ��+�D��P^3">Ң�%<�*�;��f���6ѥ����9��v�/��1ŗm�
}��Rew��q�d�[��̟���kp��8w�ף��2�{ÐWUTD�;���Ĕ^g!�m�/��1A�9�L�7�3�,GS�SY��B)a��#� "G9�\Q��>�3D�b��`^{ʜq7�]���xwIz�];��'�T��̱,��4�$nr�{C��hz�	:���0�E�>[�u;
{��	.N�ջ�x�mA�V��#K��;��@R>����#*�0��s�M�+,��� e}�|�9s[VA�R�������~~��L��ܴ%��ϟGN�~I�̒��҆%�wV�wۏ�Yg5'�TjOIC�_�8�Y̵CZ"��R{
�h�]�b�0���s�4��l	iq��a�W{���D��LJL�<���W[�xK*w$)�[���`��Q:M�he��Fj�ܢ�Z.��n��s��ֶ�mx��b,_��o�R�������Ng6C�'�a��.u x�'@p%�G��%=�%vUi=?_Yqз�+�[�%��܆�x��	�C�N�}����D	hb�#j���S烈1bW�޴�|�G�}0\[_4� ��Q���g�q��-��&/���Mp�_������M�J6��.gRmI�Bct�%�)û<Q,�!�,�̤���x�f��O�tY�\H�l	������qfِLl:}3`wek�)geZόJm	���k�ξ���ƃG�S��B�����h�=ٲ�I�"�p��,@��$t���<�up�@�)K�̋;��
��/3�A�̟M{��'���I��_�v�Y�e'?OfB;^NG�
�`���6�q�e[(&���x���`y!���-O��f��^n ��g����GPx�0�x�@��q�x��m=���_�1�J�2��6��\�mߑn5��N�nc=��5A��Ww���u���t��~Y�d��Aq��I���ؑ
q��B���V�~��؟�s��VF0$����C6C����-_���-D\����M�u^��]�Wvya~�5o����}���(�(Rc<�w��u%U� E��L�@��k�������N0`�l�Y�+/��uK]UZx������#��r��U&��C�n�V��:�-�;羀�]��$M���O�ކ'�BO��Q���V6z�x��'����\���!�A2.,�(F���=p*0ٳ��#�y��`�ZW�s5`�%G�
ؾh�ټ����?\*�|����I�+�S��l��\\��|��%��L,h"�~U�T�vҩ���g��33DWzp�1�-�nP�'��i�xn���ar��#93Q%�O�
�:�9*���%���vl�ہt��;>Զ��!����ɜ=�t�
��>���v㺃Z�K<���L=�h���9�}!�ģ��b��E@ B* :�*���8����]s�Q>�~��,h�}g�A2�Y#і��]!�ҧ�_��ʅȝſ�n��3�pei����fj}a@�$I�;	�J��hT�|�������:(�Y�۰��F��\�|f��`i�w4v�'��G-xyB�˖�a3�ے��ߝD\I��hԖӿ�d����m�!'��p�l�����֯C���H�-f*���T��\��C䘓ZSJE='i�]C	��	�9���u&�F�a��N&�TN�٣�6���Ij
�����a��5��(/��C�-�e�s!��Iꩫ�iU[&�bm*^,
\q�_%����O?i
��A��l��?tv�Sjx4h qTa�)A$�vr��l���AF�T��u暲�ed�چ�uP�����*\�:@��C�!{����V� �+�(��巻�ε�^"á�t{*g�^5�67!��Z|�g�i��^����4��$��qc���*�+ꉣ'��,�u2:�@��k`[��l�l^�Ã]y�[f]�<�h�fA��c� �3�'&Nn��#��'#ڰ�~�}���������I����
gF����������̲�,�D����?�?0�� �g�Ԋ���g����6t�y���߅54�V�	W��b%Nh�k�̛1hr��Z��++�S���Xu^灄�k������߫�	v����c�D9[�/�:@m�M�O%a[�c�8�֯��7��tL�`8Ť���.�	0J�ڼc����Xп
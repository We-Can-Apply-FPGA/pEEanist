��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@��[�nL�v�Q���<���Dxv[Gt��I����c_ypO��gE��*R&5��y�0�8l�6�hβ�r(�aI >��>������P���S�(�=]%��튇RsZ�=
�L�(����/��gx�V�e<�ٟ������'�6Wg�������&�yWhq�7L�����k����I_�Y�Vu	�e��'�u�O`�n$ ��E+=����ǔ��W~�����e�<��q�a��q܋�	�9[1��Mf��ީ����-��!�lv we�?�4����z�8�H%�n��PZN|��'ڛL?�d��O¿�l`��J�IhH�]��6!s���}w6c_����R�+XC��]��#�LM�I��@o�dZ��?g�9�Ӂ�e�+H�m�m��>i&�%�:��%m�l��J����	>D���){P�+��p��-ѵ�T�̆�K�q�u_��(Jz�\�d�=�L��w�c�B�$��v}��U������Z����Ǔ���}Ep�5kj]���x_w��>�]�%:�S���x�'��p��7J��[Q&��(��yt��ߟ� 7SZ?oе�mכ�`'P���yO���T?@o�@E����Y>�o�r�0�����?*�%`�ڐ��9�����>ʶZh���D�^� /fPsUNKw���I�k���J��*69�X�g�s;k9?]#�rU�g�H��|Ԝxeͩ�\n�	=u5�a3A_�W
��j�Y�\u�n�n��rsze��) ����qj>��Ku]�d>(�@AZ�40?KC_p�Y�O yU6Lƿ�[M<XN-|RN�@�V���b�qM: W�X�����^V|���B��=(�I��btuw
�W�Psh����,�1�FD��z�kw>g��s^ٸ�ס��mw��&[[ K�Z��o	>_^FT�O|�G%n�Ƽú��l�� ��=�3��,:��c_G�o���83�/PȤj��lʾ��!��Y�4V��f��M����A|�Mꙩ[Y�>&/��TH�p��l��L,Lr�%;6�n�b�w���797��ū�
K;|��̀_|õ��%�<����Z���"��7X_[|!���Ry�mw$
����_ۤ�9wc�>��;��J�+�e�k(�cJ�7!Gz�E�@bl>���7���+T �x(ڒ\Zz���3�*�+����"�¬N ��VôB�+�3ex�?�Z�0�b#XؽlM�R���aT�{�.������=B"�����N�����eZSo�L%L�C)�h��!h���DPZuG8� �\ �.Jz�F�A�K��U}�Z��X����m���\{"��N����ʪ�#�dɰP�FVٹlB�
C��(�1#�V�o��4�>��Q�����n�,�9���"u��uP�i�mõ��z�ٟ��7�4=��0��E�tRzwO�ݰ�}o��
�w,3{c?;X�w�7#$	CӅ��r�(�� �SQ�44�nR:8�K}^�������M���zA{�aL�����h��F�����ͫ58���Yb�,��beǨY>r`�}���,�Ɓhw�hhw�5�P��.N=��	2����E`��}�ž��RLZ)��"t[�JԊ���xRΤl�,_�JF��ߨZ'�4�� �|䀎���NQ"J(t�7"�隵�V 
������Z�5�3�2�V���zcO�nGIU�u�úb����9ZB���Y�K~Kc����X�Q���cu����F���@l����e��q5��� k�W'7zG���7��xP��}����*�g�5O�Cƽ#ol��mn�?3�pbLϏ֪���c����#Z��sx��bluu�������;���:⩭#�Wj�+v�ʨQl�� 9�s�<O��g��,�^�D�;M5d�1�D3:� D;b�^3s\ ��@Q��Nx{��Љ|�湻��A�+x�\:?�ͫ�dh�٣y=�Wsh���9V�/P�4u�$G�)2�W!������h��Z_R��z�1������bX�<╵��t�nb��^_rur�T<���S2.�k��)Nd�<x0ꖷ?+,�%�_*�xMŠ��d���P��)N�sU�����B�t��-~�v]��I(��<�`��#�
If��A��c $O�4�hQ9�s�b��7陵l����]���� X�@���-���ޖ�N5D��.���M���V�E\��}G�_��(롬N ���F%,��$= s�n!� ��[A0��AR�;_��@�������`��N�V�P�B��`��ZAѾ�e#=%����	~gN�rZ+��O�����X1��""���lކq�m�ߘV禔n��aѤ.��*�x`��.X*�s�S����D�ړM�B~35��s�M�Ƴ�{�|�#���?�!`(�"&C�T�D6���7-挜�{�� 2V�vgCS�V�-��"���e�"Z3�� ��]�$�h��d��I�%�����}dʸY����z' C�^��|��f��פ1UF���(�Pf-ĐMM�u7	Є��O"�LA�E
���}ކ���@:S¼���wWł 3���	�J�bx��rX���9We8wM��"�aSy�ʝ�e����YU/�i�$󀱚�C�1�a�mr� .���m�_+��4Th���t�#����u�3�煥��m�e������`>N�ʦE�-��mb�w��}9�TW��@T���B�\}ɔ��E���My�t�M�RS�&�{s"�t��/ZlfUy��{@$�G��@�1r+�;?8y0���E �w���$��ԭ𣏱�CĲ�J��0��X�� �Na⨹	6R���F{e��!XӪ��)����
G;�4	d�F�����Z�{���#R�B�*�ۂ+E��RӲ��9�C���S�@o+]r�q��ʫ�>��0�9�/�-L��H���rn�=�=�º)�/��T�K�\A�Ü8��5ͽVB地���.��L���0������&s#_jT�8m��{��}ຳ?�m��0f���M8�˞�����Ŕ��xU����9��y�g�&Yw�=��n�$�d�� B�b��#����M�|ދ�n1�U2ʯ0W|�u�q%X
���YE��i��˗_]�S9��|�G���R��I=KFR��Av��޹�'�:\��_
ۋ�H1Ê�Wp#��ͪE�eXUj��)��V *q�ꄜ5`�Ds?3�-#�x�=m9�bN�~��K���-zL�R6��O�.�I~�>�a�1!�Ö�h���;꡹�������Q��u�J#$�ot:���\1��"U-��n	�J-��:o�q�m$�w�F!�\��}&��++��C6�q�F�� ��Ј�.R��э��7�b�\&#s���cM�)!�$�	��y�b *�����\?%n2�r@d�:�hV?_�Z������D
�Y`��*�q-�R]k�c�j���*'������c�@��2�r���@"��(�W=_��׉V�B
uJS�fs�_�v���Q*r�����}�VZf��8��O���l��l���2�v*�}v-��ʺ��ݢA�-Ϣ�J�;(�ߑ/��W���-z�2�.`�kqYw�������e����莪9���TRÔ�/���]�>�Pl�&��ZdR�T�����c���!��,��l_���<���,�f���_(��_�Y?�sO�z$c����Ʋw�BԷErǢI.���}�Q�\I��qF�AC���'8}�J�`����@7k�:��*���M�w��=�>TjJ�!n7�}����Q?�.���t�����}��n>�7�a�$�f�?oH]/�9� $�Ho2n��<�P'����P/��e��'���6�d��'����=�r�����o��d��O����&*�bkۏ�l-ƢB�.��{/�h�1b��5!z�#)z$`eQg�l�#0e䪆�!��K��-���B�%�ԓ}�
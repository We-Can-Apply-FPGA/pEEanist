��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�8Ӝ��'�����@OI>��.Q�w2�D�봊.������D��H/X�c����ft���p��:#��'���c�ߏ�KWky�?�#m	��*`�ɦb�u�������O�ڇ��5!������mB� �C�%�#HyƬ�<R FX�x�@�g!����kU����V^�JkJW�w�/5�]��=|�%O8�Pgl� G&z�m�I���#Z�b�ujO���[ݿ�	���	���27�hP}i=�����tor[m�rL��(������t;P鬝��Z�k1�9��KN���/�d�^y��^^�lb#�c:�3}šs�M��EGK���X���n(�X��'��H��V,*,�L��'���$M�L2���f�b�9-�����g��u�~Ʒ^3Y�Sg�!��e����[���Ѽ�/��&�ǋ�i�_̰��dU���*g��F@Ѳ;`9�cV�J:���4_R'�`�K�Q1h�Ӌ^EĞ�~0�؈_Z��6и.���(8�b��I3���U�����"E#��']|�o=���m;�u�{��W�yNV& �ꦝp�/�`Z3��J���~MY�B�]�6�ԟ�5K�����m��@-�{O^��9T�D��v�"�����Cu0�'���!<�#&�VW[�L�y0>���DW9���MF�� '��u��|sO0c~|�hxP�m::}y�U51:Sr7�5�
����ZI��`\rm�L����׷i!�Ca�9{݃ofrx�%t��~l���\�r��	:�rqʀNLy�@�0���sU�����G>O7CW�7�5Gh��؜��_ �&�)�~�V��B����phȞ{�7+,�j�O��a�[��_=(����c4����h�V\Ī˃	u�!&D�#T�_��}���0�3����Ql!u�b���g.����3Y�����Kض���1��o E棦��� �l�T&���G�N\�2
H��D{���:1�ZV�}� ��M���`:>��SČ�ˣiҘ6rp������S4�2:p؜�1]xDd�`$��O*�=�s�(���
a{���^�7�Y9nàjd{bi:GĖ�������09 S �����g"cG���3<A}?�̓�r�e�r��)#^��88�t��y��B���5�]��7;�a��$�^��Ae�2���k��:���r �p��6�+�2�"����6�<��v'*;��Pk��ٵO�*U�޴F�c��rxT3�z���⬒��Ol� �ͤ<o���'��º�J>C��E��,C���tH���?Zz��i��e��T���}f��6���T�vyD��ԯ�tݑ���z���N�B*{�t�`�C�Q풎7��G��HBdC�޿��P[�y`\��"Ғ�HK�6�������-�6)+����O)�����G��3���]�y4�	���2��< �ܖ_z�-����$S^T�*���_h�:��g.aR��3�h�L��xw�Y�\��f�W"Y�#��XE��b��2�x�\|��A�r���_cm �L����Ú�@	�w��O\���9m���$z3�s�d؅Z�LW"2;B_�S1t��=�G1�+Z}88M���n�ܝpé >���m�Ф��;pm�+�Jc�׏�}�����#%������F��:,�y:���B���Bt�28m���_4������ޗ��Q�.OFh!r��	~�m�����
�͵��>!	����y#ICB[��B�k�Hh�蕼p�sNxs	� �@J��tx�F%���^&�^Yhb��t�y�Z�������8�����Цq�E�lε��{�+�5N�����o�2O_�iUj�e7����C5�ʋ�
�,���ԩ&���1�|�q��뭯mj��g��dA�[�|�q_��"�]�rs	,gw���Uj�e��RH�f�"\�"l],:,�ZQ%��[��������>�m���{M%��JB(W���[�\� �p]]�M}9R�4��n_�y�}}�g�Kw$���l�.�dTu������1�հo=�:l����rKe���UMsXr
��XaN��8��k�ױ�l�%�^1*t4L�ԙc�P�t�#��V�eq��»5-A���~|��f�hW�w1�������w4c�Z�y��|�ϛ���s���\]�r�_�U���'� �}]�H��ЈTUF+D����
䝇����Ѫ�Y��/ٹo�]Ew���t�S��i��&4���XU=$9�.�HAq�������Ĳ����6r˽�������M�QG�6�[H�>��JO��S���
�3����z��[F�ڑ��
�qOG���CS�o��r%���/] �x�ǋ�������6w�2��R��;�R8�7�8���|�~���ͳ�MSQ��`�[�)��:���Q��ϊ�/u�M$PB�o>�H��kс6����?�a&����J����G���i�&!丠`wJ�m��ۆdE�c�*���Ĺ7;��*��"˾���l�⒲���C�LS�y.��H@�#��	~�Tu8�U�e?SS��8�o��f]��w��ḟ�_��RpQ��q6%�^	���U�`���'��.����b�29��'��Gp�������Vյ�c]�LqãrL�JLp`��t��H[�\5�>3y-M��e����V[��0����/3�j������J��~�i�H1ZCP0�C���f���yF
�D�Ӑ�N�o.����C�<$Ļ�\=n����B�_.�싵_���o���O�5��AU�w��	Cb6s���gO����btѯ7�9Չ>���2�����<& ,���jiԿ�B���&114�J��y��XX^��md���_���� .�}����R]D��7��m�:R3��)��Y%2xIh`�a�ٸ��pHh ��#��JH®����g�ُ���`�k~� �D��jU��mi1j���*ܒab��8���{v�����Q�_C]��w���.J��JѐB��0��ia5r���=|!L�N��P�%���Rfv<a���u�.�!���� ����#�;����La�`���Yl�	bpΠ}��Yu(��`v��r}�"9쨇@�n�p.P�xL��FEfyPU���vv^A��4��Nf}2/��`޺�ɵ]���;��8"�s�8h9��1d\�b�#�n/����Y�����o�$���I���::�2�����������H��G���S�P[�SM.w:���<a��=���]�e�G�'����] �_�F�<uJ.�dS ��a�ꇣJNl#��?f�"��R#t�b�6״�F���Nu�y'���72��W:��ɦW����堠c��_���h�P{)�r"��a����<X�(�#� �,�v,[�+*�)��:�2�W.M�܎��Q�P3p� �oR���F?�����9�$�)7'B�eb>��b^�Ģ�FuR��nu�	����J����NuaFW�V$�y��/��l��tK�N�ثu����J��h�|m+�����»ɱbRL�cd�,�"8l��G�����w�����F� '��;�0�ײ�(R��˓�_p�hΎ!���˅��!���UY#V���r��F�RP�^D-�_��lђ\s�ґ�qH�e�D)�m����W���GJ�կO���w�)�����%
!�!�4��SRYX��g�q�h2U�]_v6��^G��q��p�b���-�ΰ�p_�.��f����.��r�26��	��yJ��d�J�7���.*�\�V����V��b:29�=�K�u5�DL�q��_s���m�Tù9
T@�c�p���0���
�8>�?�W��Z��U&���!c��s����UWt	�I=�mu,�9��[L&����g�,�l7�IQ�����~"�!�E��;�����K&�������7���Xi�t�y�����ÊG3�?+�ɪt#J���q�e������r�������P�W���vj��Gk��D��}R�
'�D*>��RGz.���Kk�ǉ�ᐣ)aّz��=G�_7Aڕ���j|0:H;�p����[9Fک���M�N/�#m�Y���m�)��M��A�@�e&ue��BK��&Jr5��&�C��#�
��e/L����v����?hG�m�Joe�[����[�ѻ��$�N�M��i\��!�ƽ������y;�CL���bB�V"p��'t �>ŀ�Y<�I(d1�Xk�R�ՙ�n�����Gq��p���m���7z�kI[ۉ.?�M�&�Ϸ���$sG����>�u������5�`�Nj�ˤ�C�x�$�&D�$��Qt q �3P��	l�n�."�k��)k9Z��:���|]2q�jsI�� %7���#��ls�09�b�z�X^Q�}���a"v �,����y[zf���)��0�`���"׭+3��b��4d�-�o�6�$���O=�Q�o���sH���FK�Ǌ��?R#cH�o<�}���T ����i��m��=�`h�8�0䠟㊻:nx���Σ�ͭ�ٽ7�L8&���'Z�i�b'�"��<��5\�1�6(���:�ќlQE����j�ȟFH��	>V/0�0 J�/��6F��=����4�>��skؒҽ�+b���U[��U������`�/�T��S�g4���g&�}��)�М�n��K	
���V��׸ž�v�6 ����\��`��o�_�)7GX_�߹-��>�S"�8�yU�6D��?o�1�� �Ȕ�`��(`{��dw*ʑh�<��V`�v�`q��U�+�__L�H���-���m���(*�N��B��4�z_��{���^޼��e��7feYQ���0�5N�x�pcE����Wz޹�E�|��=y�,�onߜf<�<˅`�zuL�H����]byw�Uq�$�D�֩�LzQ�Z��\�L�ox���+��Y�|�G�q�!�0�˧��^<��1�VM��2Sd��[���x؉!]�K;@�����tʄ��6)�H�5%4��,پ��BL>����Aș��X����_w���N�,�`�4$�R�?��f�۳t�I�)�8�⇂/��̫��*0�B����x�@�	Z1I,�%�H7�Č(��Âߪ1����;Q�t9�HU��m���>e�^��<��wΚ�& F+P�.�eN��Ѵ�~���� j�����w� sMf����86���/ˌ�HJ�I2)��r�Ôo�)kfO��&�<��r�!Ij_g2[/sY��gU���Em��X�7�R���`��*��v0���݄*�{G��=òQ,�\��k�>;��a�U����Ą�Ǡ��m�z��h!��	]�5�1�A�^�8�OӶ�5�����F��$�#�Սf�5֟�{�^;i':F�[�I;jԕ�/�Ag��7�Xi�����9�����`�2P�ZT������A7:kG�Xs�$�]�mw�8�-�a)>#೼���)3?[�IX�MEa�,�?��2tJ�-�d�K���(u`����߂�@���j�k��#����D#�S��=���q�$)t�0���T��vIM4��fRVA���>N»*4��	_"L��2�·8કxO���(&�[�=�"y���@>/[w��AQ�8X'�4y�~崛��=��r��}��)��F���a7�քe �)%}k��-����E�����p�G��
��X�'Fpm���o��YP�4�80�B�~㘡iG`{d ���c��3��@��1_��0�с�렙p���c�^
3��36��I�"������!	H���y��RyF�T�-J{���K�Ԍ~Y���oy�8�3���U7���zlw� ��;iHo��j�Jv~o�
���A0
@M���  �_�a�A9�x$v[J�,�Ѳ�v`Nd.��<�.m���k�W�������de�2`��B��1$ǭ'��>B��Й�|�VE�����r{tɽ������5~2��1�m���al�mJ�P�4��ѐk��>���ic�����˔}b#-���a��Z�� ?'3�4V�0i��nT��-�0�mM��!�ˆ�[HNAgͫ��@���Z��v�9��=t���I�"C��� ����Jz9��A��k���G5*�o_l�"��&�a����3W���B'��g*vƬ�m�H T��:PH�3�̕����4H(���~}=�tb(t:���i��O$��v��b�t��X���� �[E�y�l�Ҧ~}�IO  �n�sÀ���Xk���z0aN$�g�#�M���l����B���Ux\�.+q��,�g=A�J�?+�췤s�#ỳ�^T⩘�VV�}�i3�+�V�a���Jrã9�b�wFBX�m+��V"��{qZcYȝm�lƊ��v�T�PEW���٨�d������I��-�S}d0���7�u+ ��J|�aK�.N!aР/����(�_3�ms3=@�x��z�pB����0<����/���]��i�;�2E×%�5=���Czۿ�Aۥ;xP��>�߭���'˯D��'W�q8ڻ(���m7?������7�Y�I7R*{��H~��o\H��#T�`�})Os�kqO�#c�Nk`(�YTy�?��h����:�8��x�k_r|��*,8��Ե�}���^��uo�w��"zu������I�{�W�x[6v�h�z���<�3�T��(CѪ�>h��)=Y�d�rɘugH��ׇ�۬���yA�ޅI5��}(� A*�-�JPC~y�7O-ԅ����yi.Y���Y�	ML�(��%�C��e_s^�#T�5)�I�f����9��}���\��y}�]�F�,I�_��P��W�z�R����8�}�<�.j���큜;rP�WQ��Ґ6����kr��đ�=U������X����<'��af���N�í���,�i��B!r��y��
f��3(Bu�9yk!�6h٘�f�9���-a`7(1JW��Xo����Î�]�M<f�*�E��y�q�Y�m*h'^�E������}@��]K��9tf6#���u!
���	�ݽ�\�l� A��C}�6Y"�U5~�*�P�_�]|E>$�O`B�$��T�{7L7�tWl��)Iȝvb���4S"����TS+2�ב.�� �g���Ҡ�w�^N�P�1� :�'�,f&>wT޾���3���g��X� ��$�6-�ՠu��}�l^�<��l����LE�W�]��r�Vz���S�˂�ٖP��(fK}���'��g�?��ބ<��&�t��3
�b�M�c���й��~�.����ѧx9��̫�r?��4�������w�_Yk�傍����qB�Tn�Z/�>*��Ȗ�'/���!%G���k��C$T���U��*&� U���������1�s���fY�����p��ɂ��~ײ������܁�Wl��0'[�@��i^ɇ�D6~c�t��N��z�8�@-���� ��L̮n	��#ȯ.��a�����x`<�\�
wV>g���ɽ7*eP��#�8Q�[1�!��C�z&���Z�)� :�|(ą������}'<���]��6�s�yp�bvs�ܶ	W9W�H7��F�
B,'hD�ہ@
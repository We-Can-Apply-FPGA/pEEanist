��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�t�!9/�f�=b�:O����}q#�����ʎpH\Ju���#y9?� �y}��8�6<b�5-�l���Y)|A8��'��|sx�����g� �
�N� ٺ�R���L��0��eHXׅE�M��7��o�hMj|O{�	���{{C�J���L˂8D'�Ʌ����%t��z?k�.�l�]�'�'^���_ч��w�(���[g�+���V��6)�gc*�^�`<]w���M���7!���rZF�^U�"f��ď�
d� �l���V
�uS�;���n6�h �S����P�}3{$�=��}�������:��KX�23(��ӎdMm:.JN�����|��G���p���mQ��jL��N��ҙ��CB<��1�H�&�Z�lC�Z��k4�u�7�? 0�$e�x��j#�:�4<iO�������|a��p��a,�>	_��i;2)p/�4cā����(3�
$���2S�8=��%#��YNƜA����	A�g ���(Bf��1�^�F��էIډH��Y�=��pI�&8���� �2M���4�m��C�,�����=5�!�}�$��A	GX�W��8�G�'cQ�g~EQ�\��O�zvBR��.�炁P4-�Oj���M��e�)�ů��10�E������%|�@7T6�,+Z��`����=2���&ђS6�R{�2�s�e��H�j�du��WB�3�-!AH�'��=g�.[�|�x�E$�Z00���Y�4�]W���	�?ٖ��F�f�#R�9.p��RE�4��� ��ajQF�A+Y;�0'T�Ы@j�eO��+�Ϳڟh����3�Ѣ�K��P��1'M�W�I�t��E�V�o~H�un�n,%xYS���#�h�ֈ��.۝`�� ������XE=w����-3��Ţ���u��w�y�D�
�*�2c�7�#�f2c����װ�������f�zUs��?.s-��L����hPUT��/[X�>������a��EA��F)����Jͨsj;90�YAs�n���A�i��������xE�H�%l��`���Ֆ�
Y�,R����(uUQP]�Ng*#��C�ԧ7���G-�� |��]�#�އ�h�|�{*�۰r�����v�}���䎧/�p&@o!����P���W�5F��"z�����m���a�f��t�#w��F�j�՝�Q��	�u�l]WM֒b�vB8ݴ��mr���m~���z��A�i'.���D4�}~ 8�$!��[tI6-�ߪAm��pя4	�	��_RiG���oe��/z�s�7]�M;�4v�o��!�5�Y�Q��¹���	�@�%-3�]Q�A!����e�d�GFF�E���n��IW6.���ь�TqPG4�
(��/n�8��F0�pP�tG,�+ �b�b�A��y�hl(�#a�)-�^�ټBltn�9�I�z~��������)��حc�E��W\T��ӫI���`Z@�=��h=�O,6~Qz�Q��_��۞�r���B�\�[i}��k']���g�fQ|7�y�2��n���J�0 1��w�}oo��/*C>�I�=o���90��m.&IP�H���Y7�)�ȣ������,���/��W)�[d	��J�ɒ5y6�(�~��+�ļ:��6z�)!-��G�G���ӌ4�?O�g%��F���T&�p��s/�=D��=]�Fe��o�y���D�"�酀���?pim%��N�Q�j��}���U;��F̉���n����AT���!������oM�S<�-C�%/�!_fߘ�ٺ~z��eE�h��r��Fk�op9АWU�a���c�Bۆ���7�#��p��#��881Q�mZ�!��j\�?
S��K�S7n�9�*���_Sr��'��d�ۥA�9�����7cW����ubY�RĊtUv%����3#� GE��T�`�J��dLn���9S�� �א�\$�2y��+�>�o���g��8���� ����у���j<�~�(D���m⮺˛#gѥ����]���!	Ng�4�##D�Z�蛮�m��@6������8����H������޼�6�9��0�Z3��;BN�n^r�ÎͰ���^��N9f@y�l�xz��ȁq��}���e/�K�J�%gf\�)�6b^D:Y(<�Q˅��0 |���vj±�G9ޭ`�D����T���� ��K�&Е�K��آq�f����3��6�?5����Z�n�� ���9C`��06Cj��׷���({�Q�z��(�	�(5e�c��-������!�_��rx����V�;��H���j��1ٓ��J�������O!�]F1���|5�q������^/`5f@XCgcck+���*�Q�uf�-��+���Ũ����a�K�j>Gt����M�h�lS�l)��3d*m�7��!4�
�2xXtO����j^2U�X����Γ�� �8v��E1��L��1:�BL���u����1]��c�q����u1�6�Q�6���IU��(ـ�
���Z�Iw�a��$v׿�Y8��AC)~2��ʔb�0N�n�� iDH=ۘqN�s�|E�� �x0��V�ނ@��au^�)�er�Y�$ASO�MC�~D_��f��璮�(��{k/������B!R[ˣ�Y��'ߑ>��,��t�b�:8&3LY�q�yv�m��[���F���y�}H����[�;ɺ'�4I��B�΄A$y�∐j[����G�W��ߡ�8s��LX;ˢF<@Я6W�Pػ ��y��l�����l���d�(qg��"��]&�7�ϥ;7��0i�r����W�}}G$%t(|j	�<�������J���:�t��㧹 ����)��Nv�ũ�0E�IMS.�'Kt|�y\WK�C| n�:e��-*��*�j!���~�h�_�Ǟ X�L҈��'jAl;ê�h鄸s��V9sXc��_'�SD�ٯ�1�$�������:F�;��5;f��Q_�Z�cKA��$^hj'�D��F���b�6�@������� ��G�Ʀ�QD��ް����\kF��γRT�5��b57,�mjo�ˀ�'�}�y+�A��� @e4��t��^� )�(%�C�\��0fλ6��_V���f�%Q�jL�R*PM�����>O�����C���fK	�F��du0]���T�tI���U3��.�1S�[�Jİ<*��F�}�T�
���ĀA  ��t��eH�ֺ|�_���hj�w�xN���`�:[��|�0_O���������{:�.�c��6�U�U�}q�?Z�Xݏ�R5��Y�Ë�2�fF�%;W�ͩL��Cb��S{�.�~ܧ�x�g''T��پ^а�'Bg�\�^R�+���!
�TebMbbg.&�H�z��u�'�=a^̱���L� �W�Z�7F�691Dܛ������v9���ɢ@����$8I���j#���%;���K��S�HY����ކ��x�G�M�n�Ǵ�UBؒ�2Ұ#ɶ���)�61b�;�F7X��j7d"����Ϟ�ҲŷV]�fG�1��7�MM�3�&y�9�<��y��d?_�?�֘V��q���ֽ}�цh��ʅ���j/�~�x_����)˱��������!�m��)�H��#Dp�TZ�r�f�vt�H-�� [�  �.�>���W�p�tT�j=|�YѠ�k��fit)��3���L�O����#�[��+��"��-}�����Q�LS��Ҹ�@��:��qPC��G�3=M5R�;>�}�%V�x�eޟ����u���L'�4Z��(/ᅻ@��,
�L(����=�|iQ���9S4_N�ܩb�.��Ǻ`6v�r��c��!gFy��zY��ʋ�-B÷��	�ܐ�{%�~&�gT�8ꖔu��y���8qa.7#���Gڒ����@�:z=�Z�k�@�L���3��	�Q�pl6n���%��_������e+s��}��y�@�� o��̉<ڠ����K!�-�JE�S2=�����Oxӥt!�p�z�ڣ��b���A�[J�h%��ˍ!�!��[����;V?ǍHt�j��Յ��)��!s�u`9��Z1��_j�_ l�8�*�3�Yhq����C���DN}m����a�,�2�4�د�L��.��Ӟ������/�h̟�26��v�2K�5����/��L���(&T� GN����YGt�V-��;e �W�1,-&[�����, �%h��b���Ľvܸ��G�@�gL����
��>���������l�B���9 /m��o�*{ü��!4xc��y������31J~��^��x  HH�Oo�(��S�uZ+~��}���ʆ�������3(�L{����uqi:��x8�GD�t�°���䉵C�D�t7Yq�1� �3e'K].��e	l2�U&;d�>���p�eQ"���S������|��=Cm�`���҈Dn	�J�"��2��a����׎�?|
��*7��2/��N<Օ����[�.<�1������T�׺�Ǩ>�.m~�^�a]5����W`4ȧ�$�����;���`�O�� Z49��ɾxq�~��x����q�:����)Z���.�Ӽ@�RI�ިM���6Qh�y<�;��d̐h���-#�R ���-	����&�a�;��&qk�"&���U�4��}�I8�>>�������"$r플��y��'��¢#�EFI�ڽ
�ج��W<�=&�����!L{	��S�n	v��'f{��{�U��cw�3n�d#�����D(��>4ݕ�K�מE���d�D�1���|\�X�`�+C�ў�}�p'9Kg�0���~��J���� \�O���G]�w�J��W.���̏��a���qk���+��L��Xoc���<p߲�C��1�.?^a�J���;�`ĭ�4��C����QQ�2 �7���s�� ��*��tu�
km� ��O�TW'C
�qT%pC�U��*
����e�M�4��	�S�ѓ��`�m��m����Oܓ�{Se~��T�Ie�>����~��~���CvC	�����n����o��R���J4h^Ͷ����ץV�����t�)@���nʌ�,�K��'-��jY��="2Zx�`U墅M+�GNt����o�,��h_R�J��и���t�IJ{�z���ml��#G�ok�8r4+־�e&P�M��f��Nz(K92�|gr/L���i{Sc;�Z�2TK}��U4�#�p;�9�fi����*�5�/���Ľ�V`�����W�3n�ʊ�	��G��\�%�,g�홙9�
3��h�o+��Mvg�`t�}����h��F�ll�59n����忺u|�j�Br����� nH�\ɤך�����ġ��fx�F3�$�St�[�?rO����r��QdF����M�����[�d�o���u��|?D��g�a���ǸjR�\���@��`b4uL��*�O����i�3�0f+m�}4�J�.��EU8'��q�yR!��;�c�n����݈Et� ��i0Yt�u����B�/��f�L�V��E�>j�����ƭF�@���2A�����C��D|��}��v ���(�_U& ��]���P*�ټK�4BR.�a0E���&����$�@�M�:���йz�/���wZ.�
r;�����(�.������ku/?��U�2���-�
c����y��|�-^���?@ac���4�>���r{W�>Tj��p.Ҿ� =�ށg�������- �,���(�q�d"Ł[8���x�{4��cJ�JQ		��z���xA[���L4��鬙o#�K6+��**�^I.;27�����=�#X�":+�T���;"�QL���~ I��x9�}���)�a���4 �ɔ_�Ʀ�Y���,��z��� � ��o����N�M��j���P�~���=E���&8��a˘	���	�Å�Y���;'N3�����}F���f�A��:��~�4��ҚV��z���i��U��Qz��U�5v.΃+D1��q`+	�Ѡ�����G+�mܢ	0��3��H+�ΤV^�����w����5�D����~O76�ݺ���v�<��y�m�~=Qn�1�]P�r��>|�#��e�l����`
�Y[�LY�a&L*2`�$=����N�Y�4d�<��K����Ի���������#Q��|V�W˟�m
�g�;�UsyG��I����Z�(w�Ʋ��l.l8�_�����w�:��J�ܞ �o.��ܤ����R �]Շꪋ��F⻆�κmI]�Ջ�粣�z
D�Va�A̐�b2;�e��i�Z��'�bH�K [V�ŀ�����;\�Ά�qv�l��t�ںW�P>�^��W�g;<��%E��n�$e�'��]��g���Q��g�V1��@�~�|�ɔaM��xbYqm��[�<����� ����2��ߩ�Pn�$^�I򐘵��wh�K�'r\vۚ�/��却�r�$,)~f"��]���(Q(��R�w@�j�׏����)��f1߶qjT��=��* 3�^�gbf�j��(o�NE��k�j�;���_8�*�q/�sxao� �0t2X'YjaY��ᨻ�?���^� �K5>�rˏH��:*�c�M ��T�eq!E�t�j�����' أ�H�,Jʍ��˹����2��e�9��<���KQ���5�vBC�RfӤ>�M�����X�B�O `�[�zc���j ���@{^4���g�gE>l����~�����N�<�mkZ�f�q����!��h��,	����~U�/;ƍ5�V�� ��BK���V��	�5�7��@��$/�/A^��� >K�4BM}Y���Q71���|��K�d.�O��2��}�Z������ds&���E��{��]��K=<�����'1$\��i2GR��;�Dx�R�	 ���6�f��Tؗ X图#y|�,�:�'���]�'�#O�H��%r(�~-���r,�c�i,r��\�t!c�?E��v}��W�>���Ot��^������%ܥ�ai�H�3�P��џ)�nt��zݲ���M���_�v��	fT��x=�j��¤����YI�	�Fa�J��@�O"�Ɣ.x��H��~[��l�p�;���B�2�{��r *�9�����/i�l-<~�}"f��k5>ƭ�g���{��P�5�{~5nA�>�z��j�;���P�/j���c����^�����TR��;z�M$�}|���x������
E#�Z,�J0�U��?T��ލ` ;`*�zw)u|l�"f���:n;�{Ȧ�W���� |]g�p�0U��:�󱕙��B��@��0�gq��V��_���hb�f�#�`"V�&8�G�C��W��_�*W��#Z�H7�3:O�tҺ� c�̳�46$��{������x�X-7t�!-W�f0���/�q��녧�A�u^��#����Ѣ�9�M�=
�1j�L�d�˛!a�.�1 *�6^�x�NԔ/B��C��G����_��m4ǂ���`�jv[��ޗ����D�~�H)��C�P����$�/��w����c��*��⪒��V�T�%e9G�<�)��#?��|����7�jmߚo\?�G���R��.�����*��5�S���]4�%�]�5����g_V`���K���B��8��Z�A�D�\��MH-S�&����̤`#��@���ũ9��ۿ��-/�A{��R�I	�w1ѽcĐO������Ҟ�U��F����&���[��36f4L��`�oj���!�9S��7I��ӓ��F;G�"\<HڼF���h�XtHn���\���s���F>�=4��W|����b=ߙՉ�YŢ^�	X	d��6��6�׺�\��ȕ�sC�H�kX_+3Zxi[
��.ucs��#	�c�(�wq�@�1������y�nϝ@����*��^j��Ow��/��V8����
C�(y2!��!�bo3�/��X�=�t0�"���%z���aM_8�db$�R�TE �箲�,{�A�E����p�0;�� �v���ܠ8MT�Id$9+��)���um�W���H��+������C��5S�/
f�YQ8M��)��M7�\����%��)x�jo�,��E�4ؙ4��}���\�(ݞ��z��۾�X�J��Sl!^�x���2ܪv����p`p�Q{�4S��n
	Ѧ���iy�ӆ��|LYs��*o8V������⩉5UP/q��»��Vw����8@n�n�cFTbx�6��:�B���֮kh�e�ֳr��4�ߙ'�*�c6X�)�T���s 6O_��,�[�7�8�' �R#���l�%ލq>2�_��D�,��A���\������g!v�F��%�W�m_��b���>�'@	a�����E>��)+���R�}� ��������.eKV"Ĕh{�_�y��81�z'<�i1�����i2^'�|Y=b�ٵ�$�Q��μ}R��H�Yd�-@�%T���N��}�k���kʞ_q��.$����z�ԕ������L����@b��|��a�Vɘ���1z�K&���3��T�'��M�A�P'	� *�AVIm��k����b����w�C�£u�WW 
f�>�����20's�(�2�'�#P�Î$;�s��uf�x�9����#\��<���E0�9l�z��'�3&���y&�L����͇lf@>)��y�	 K�����g�ST��ɸI�]dѠ�����})�!+oˬ�=B,�-��$#��<g�p�����Q+y��ΰ ��;ڲ�m���B|��My�m���{S0�E}H����Y�Vvdl��J=�|���s�H��F7�$��$��P��r:̶o����P���L���#u����M��o]Xծ���{�pz3���S���p=7� �Z$UZ��`��˚ՠK��A��iU�/g� <ƌm��������W�T���?�$������V��,�'�ۭk�`	tHR���v���x ׊��x��J�{�V����|k�/N8�"�˶-3X�,U�(������壶��\��nͶ����I�x�o����:Pp�7���ᐛ�#v߲��N���a_�+?���p�ū�@j�8�����[S1�}X������_�0�႔��v��ɼ�}HO(�4T:�Ji�3! z9�y�fkB(� ����ɶ����� 4��<��(3c�1r��g�Zw�|Ų	9�(Ӌ�)kC��Ҭ������'oVM�z�0�E��+�G�i�a����]fج�Y�0N��`eű�g��4�i��0ojKZս`��ɂeT,F*�?"¯���������]�z�Q�)yЗ�Xe���( X$:b	$Gg���b��Z0����X�����|;#R�����Q�ﳡ��ˇ�d�߶��I�~��%u9N�J�[�$��R9����iÀ��I�VE�a�3l�Ug؇$�[��q`��??�I)Q	�� �gm��恂mt?�|B�/QN[9���8]"���Ai��VM�*S�8 �9k^��`aG��%ŉ���+u@9�^w늉v���Y坁uF%�=�B�tzC]�@?H#�f.��V�.�<_W͸ĕ�I�|ڗ��'���K�󣍽Gw����q����NT~,� l�/'�7���rS�7&���'�)���u� |Itݚ3d-�%����bR�P-����u!��,Ce6�:?�y��mu�~�L���`bE�e��i��7]�\rF,%�ʲw1��)�$�W4��R&ف�Bm*(j`��I(�~�T>��7��Bmb��$�q!�We��?2�4+)�?g�;�ynA9!�GK�����  2�q�z��w��u�_sX1��4&�b��3�V��I*�^��ކ�áLR�� ���[	�|$�;f.�ZV�H���ک؅"K'������c<h�+u��{��9A����xC��T�d��+������ί2l���#.��M[fnrt�T�cC��ѴXus�q難�k�T�TVg���}����<>�:���D}�pcv8�}p�Af����4t+l^�+��)6�����L�m=5��7f��.����)	�&��U���fl���;�n����g�6U���]���͎�D��oS�J�נ� �!�{��b
W&���,�����B�Y����թQ��Յ��Ҵ���NQ��ܬx�dDhi�pF	����j�s��~���9�σ��� ��>\�.��;��� `� �Au*ߚ�51Ě��G�k��	ڨ7�7\I�߼&�]��z0�͸E�FL�F_��x�����?'�(� �:��TG�rڋ�Zc�%i-�ع,��d`ڧ��K�����)���/�ĊOi�Q$���f�Q�ᄰ�e'�<&/��s��$���9�2��:I��"�U͠�I`����n�5�1><��Gk\�C�9�KHq�{I�Ϊ�2�.������2�����+�qIKؽ֫���/jJ�#�;#�[��;YD!*|�&�I/�D�c�Yo�6�0�����D➎����K�gglU-���)��4@�D�eP�&!�p:�)�B�����X�ߨS��1&5�t�f���I��ɏJ�2�,�`?�*x���銳s㝦�%��V� Z5|y�D��p!��zRp�c�1eS��/Õ�;o'��%j�D���-��vd�;Ge���V^�Z�4w�3kh>p��0���N8"�:W�^Lw��tg!a}�a30j�t�\l񳍓��f��0j�;���j�^k�L�����5����A���5�	�CH_�k>�P݃9!�6(�j߶��E�U�Lt*��	�>�-��!�EV��ޣb���2�.��N,��#7/��{9�%4�S�]�o�]�m����	��'���R�E+_�(�,?TNL���k5qL}A�r��̛Z�R�3v�e�L��'�ȵ�a4iR7l'x��A�ڸו3�g�G6��o�B T�������q���N��qZg��;��(dxK��0B�m�pH�#cv�X[ܸ�2�AEj2iT=��Q��ҹ��]�l�*r����+k�Q ^�m^M�[P����G.�:1��R|��� 9$=�M�������ŧ7�E��	C�f
{ʩ�p�L�u@��13�K�jV��hn9��?����e����X!�� ��|5"
����6.m$������
(�/Z�4i��lb�\�4y�-��%�SO�����{�.ˈD����6��Lɡ!P���> �Ñ?�L7T"�*AcJQ�*���,��afj`۽:�9���;iM����w����G?���č���`k�}���i>wuX$�cC�z�wa�7G���8���
�.����`s�a��������|u�f�[���C��4R��2fq�)��5��P�)}��6P�
�����BA�,L�Ts}��Юw�b��%�%m�l�<)�Ù�����5	)�4[JV!Ig;�p��58�F��$B�Sx�cj��m��lOEZ/+,
�N�}S�ʒbͤ�W�=H�S6Z�{��X*d��Tݕ$nH�90;$���m��Q��������`�"+�+��z��QZoA��9��u���	�8k�zG�iY�)���a��2��@�rj��x�W��Q)��B�K�X����N�f�����x?^�X�O�=W��,-��8�2�G�������nϷ��V�yK�^"1B1�Oв���D�@>���K��1Y�u���Z��Ѹ�B��\�I�@sN�q�엔��j�����@W�R��g�stISn#�䜰�&t ��]:oǊu[��_�W�������� �������o�&�\W�|��^y��W���Q;s$�
�
1����$T��l"��#�t���t�=��]�w�.�����%����V~)r3VJ���y_Aكr�n&�WbS���Vˊ�wf�pD$fN�b0*~Îݢ���g���.�<�@��Nd����dؚD9�D����i��y�~$���Q��s�[JmWc����DS���A�"v4�=�v,o�)4�:�f[sd�n��I���fU�p��"ݰ�'���"��;�m%�v��]�\��y>H�j�f�W��` =O�-j�.��'�~��贆���џ�WE����gX~2�{���`L���XY8T��r;��Vѥ�e��ryc�D(����`Tl���R����f���ħ�ڜ37�Ս�tv�nB+�S�j2��ص5������4�V>eȔ7`,Cz��A��xc�1����u,2�/L��5>(�R�<�-9;���+q��M>�*�a�#������1����.2������֬��ob��E���k�F��\������I�g���V�:��Q��;^����,�/=��=�>�*6+Ԏ�?�6:<K��r�;1 jc���,�f'/9D�a��!S�&T��%����׼,<��6(�7���y�'�#.fF�����Y��B,E�tù�Q}��;���lF
=Ri1M&�9[dQ�ǂ �ˎ�0���Mwc%�����Zg����� �Wy���~A�%�i����&��#KqQM�GV��hEN�-����!��A�/��t�oy��o|�R33F�i�[������7ؠ�g"_-a���N�6�$ �Z��u��I�aÀ�"PL�4�o���KS"aH}BK���i�I���X&h91v�@$\P��?r_pa��c�����pLj΋��|F�K9�@�VӺSp��q�n�vFq#K� �э�d�P�� ��I^�OD����)}1�ܖ	ҩ*A�̯ZД�q��,�WÃ��fA�Ez�{��b��#��x{Q+��QT��ۈi�hL@jo��l��8u�Kg9"C��De�u��������������Wp�jWk�3�~�7Bң�:Ei9t���W��ܡ@}�k`r]�bQ�*6�9����o�Q�#ְ��.{N�W<,7�p΢��=b��7��.�2��92�$��Y		ٔ��4b��"H�u���澈&]d�ae	�+V����Ӓ��2_��YN�h<���TN�Z�Ӂ����m���-�Ď?B�W�D=�'�/<M�KFПA��&�[k��1���K�j�!Ȗd�Z�'��e����;N��@g����D��"�d| D�M��^�1 ��8����������)�Y�{��[�KKi���U��]=��	/������]EL���f �i���)�%pva�pˌ�ƴb	 �5[��"�f�o4i}��.�V`��a6�%�6ԅw��}?6�����?u��j>�-�U]��.��v���s����&��Ԯ�z��W��W�۔�c*&'4�~<�0۴�Hop��%0��Hq's)�d�����C���f��ũ�Q�+��0p���P�.-���aZ6cTN�Β�}:?,�둾;�bv��{��,�7�DX�x��o��XR�٢>���I�xR��l���{�ڔ�".���Jo&�Fڲ�����!H�-.�������TB�R:��z�w.t�����d��ah��0�yaϏ����Q�*�Z:�bgz���D�����	XP�3} ��Y!U��cN_�%�W{hе��$=7�N+��cD*��9�
��ջ�"G�Wv���������_o������`H��*�
wn����+a���\�^��|):S�@B8o:6�n��}��0%ʩC&E�EQY���'��ZA��˗z��n��ʡ�zn43�~q�4L�;K�R�p��ef�D�0b�b̑2}Cݱ'%C4�������}&2b��0Lp&����4l��\�q=?���
�n��f�O�*� 0&D�|��u	~}#u��`~��U�"u ��+����0��@�t�җ���(F�b��,:E	�b�ݢi&�[Y������M�^	<����xA�I�O*o,��0MbFZ0�V0ף:aT�'�VkC�c}��1A���)K�ϫC��]{w����A�'aPܘK�	^*���۽����O$l��6>���n2��:�b\S��J�Ȱ,�\����?�d%IO�j����qhguTS�R���*e�JS��I\��/{��U������>��e��}������@�Ʒ��3״�\�f�!�0���N��������,�lF�t�V��J�o�k�ef
#�;�l"���?�M��s`�>����=-�w���ODԇ��%��z
Qmvb�]��<'����N�"<�! I
<K���� ��
o����ߠw��#g����~�d�¦EZC��9m�ɩ���q�٧��W��#�3�o�C��3_H�m��,�(B`f�Hp��k���4�V>rhh�K�^Ha��
^���B�_�~݇h��	�@�V�zLSG�'9-�Wj^5��	�~T:�?�}C��8��I��F�P���<�f�)��ٱ�v�9����Bz�ʥ�y
1�aG5�H:@dp �U�Ͼ �a��2&����ϝ
�����i-
.�az`t
Q�\�b룧��@�h�R\;�Dx��j�KpK~tM��	���1�DIG�};�<�����\�k
Dܐv���U�h}�C�5�=��R�q��ӧ�{ʚ��Zs�pt#e+��ْNOo��@�ϱxZ{ȳҼ3B �8�i�G40��Bҏf1�nB,S���u��.�{*"Xߩx�`e^
�^SST�2� �a��6�n�M��~?XRl,�3�WU99�ራ��I�񂅴�ʵ�,V����5�g��,D
#|r�D�y��Y}59�A�᭚߁R��#y��R�pYp�4��ڪN�D@k^b�I%?��?bP:��e���I�ӡHP����5V�=7K:�#H`���]gD�cI��.ƻM�=��9�Ž�j��ш O�t���>S�S�!?{��5s�<;�#�ˋ�$,˒p'�R�N�9Y�v��q�|�(�yD	R`���	!%G���XF�����7��K�T���P�����@f%������иm��Oc$W�y��,s1)��ZC�`@�ю�P$D\Ԙ�+�ΊA���&�N@9�C�冷�Y1��0J��i&��F�>��D}�Ò�yR
�ؤ���k�(1��������3R���W�R�p�ߧ��ɭh01�ղyd6��G����WQ�2z��$q����o
�`౩g�'���=|��{Ԫ��+"���wH4DLe�H����]'8�T<�uGK�.��H/6����q�E��M�a����Ҙ�&C�����Z�TKeH�7��/�h���
c�j��ˋJ�JL��e��|X���e{��H�8з[=OYR(��6�V%p��Pw;��3��G����>�kN\�&�fYZR��Y�P(��z��*i~Ok����9�����*�]o�f ��tKj�v�Tr�QY�F�^ڗ�*� [�̮�ޫM�/�
����LZ��jF�-��J�$��÷RL��\����H6u;Z���vt�̧��غ�W^�T�xC�%����4�?�,]4����^���ڗ�%+�Եٟ�L�f.L��x����N��B���1+N�qC�M!�V���n�F�b���>Řaӎ�����ʳ1D���M���9�'a���.�xtH��-�W��p�Q��lY��S�=}�N�L'y*@�����V��[��ں@::{����m�r��~ۨ�{Zt ӂ���t39��=7�o5���}����c�ʯ�ڋ@w�ǆ�6d�#�⏳F���k��ʄe�͝V��6��M�L�ܑ޼^�P�g�E���d�)5�&�����U����٩]\�Pw|A_�I?��cr��a�ܼџ��^��7:᝶�2�3���1��a�V�-:"�&��Cy`��/��FIYi5R�j:K�8�i������@U�E��"XiϬ�$������/>�6g+$�+�1\$O�H'ߴ�^Q�ȣ���S���ٵ^'6E��8'S����6H��G����r���Z�e1��m0�@m��d����z���!� "�ӷ䪽�q6�������g�g(t�#Q;L\��C6ݭR�;o���b�! A���Z���4���S����r�Z5qN����x��4Kյ����I���+ts9�i�7QE��{:�0���N�h�q_�\X���k�9�
�6�^�Fb��.b�)��������6:fc��;n@�0��5��.M.á�?Vٜ��B.�9)E5ݝ����~��촱l�n�\���r��15��@v�x���Y�+��t9\ab��9FI�QՖ�%�τOײL�nsi�O�a�	�fx�W��_���V�N�C�TX%�8L���"��Tyo@�(�T,��=w��B���n�x� ��w�c�U�AHV�dA<�޻�-z��V̵�<�N���X��>�}*~��.n(S��=�����,��^WڀyO���]+����+w3�1��g��e\�����!\�ڤ�t�QZ����O�|(��Ōd��_�O>��sc�I,;�S?�},w��w� H=��V����R��6Vļ�jwl#/��P�J-5P�4��()�d(�ͫ��c����:��t�L�3���Z �]_��Ƹ���C��SW��<*��0�5={�*���Cx�ȳb��H�$�i�K������ߩ�`�>�����|��/)y{����tU,�C2�1Ի� �\�6��m���O^��a�=���X-,2*<~Wڂƶf��VT��z�Nӿ��^�;�	&�0B5��Ф���^4��Z;m�c�+���sYH�By�yOR$�_z�%m;�N):P5V.���v�#��Ӕ F3��7T�Ԇ�H���V��>������<3_�|p�6p���P��	��ٸS���+9yv���ܰu~�7���=��F�Q��/h�ne| �O�m��c���JwˣE,�N���A/7se�B9z�|�,��.KQ��#x��:��PcS��m9�dѲ��.�3x�lU;�'���>?�A}	C�����->D��4*���3��0t9!
��^,�2��	�dv����PW�Ί�f��wd�@��R��M��?*ь�7	g���*;u��r�Z�9��������P�ա6y���܌_��O���?_���'kc��������k;)�RܙQ��p�Z�/���p5�o�Ui�6�~��e�	�iߛ?��zu�P Ƣ^��4=Ac'�)a��-����o ����p��P'���0�69[|i{�Ԇ��9gs���8l��G���=2�Χ?��*/��ԃ3K�?`�뽉(`��cgܧ��(hںԭ���鱼���r��<pM��u{�R+��Vʨ�"_4��C�n�׭�T�3'Y�X蕞�������(�z{1;=�}�[-i��6y��v��o;)����9��i��@��ݪJ濿��1+�f�/;!�T!����ӌ�Yڄ���V�����;�9.�YV'��h)8wt%����`����d�֑ɜg�+�g�J��JBc�h0��s��0��������Ƃ��\_��l���ֽBV�/�G|�VM���~;(>�tƳ�>�L�{���Y���ctH$!X>ʋ�pϕ��ې�w�Q\m�{���n 7X���pW=�<�r�u�N�'<~�Rw
�D�m���ې�%H�=V�^����Q�5�Bcq̃$4\�/�&�$0>8�b�	�������2��4]ne�4;�KgXH*�DP�� !�I*j�����[�>�;m����B��1�U7��1�㮴��9��i븺>��sH��CP�L_IF��p� av����>c���Y+b�_o�F��m�ޓ��e�7�-�11`|K�wi�6�������7��[��%�����S����x´ɽ�[������%��kM<�E(l̵��@k*�:���/�*JB�*����̺�Zp2����=RI� `{�����oQꛏ�������q���惯���2]H��=f����{�5�,��l})-��9��M^2@]E;����)���i�عY��&)�T5��I���J#��h(�G	�� �����#)�U92����H�%�����8r@t���l����Ű�~H�)g,ξk��a.������
‍�m���0+���|$gSZ�I��Ko�ĢjGy̵yV��ō��������v�pr�	,�U���X�=.������ۡ�k*8��ƛt����J;�ih�g57�=����=��T�4BVmOl���*�2�/�=����^-e��t��6��%h��(��4fL�X�0��3��A�,��3Q���3X�?���Z��q��ga��\ʦh�NyX���L�2�ޘz'��-)��%�NG���0�0����5�7��Y�qnV��6I'�k����{Ӓ��%P�|��5f�B��Hw�n��?���H8��%n�@�p��`���{k��skT��&��i�D�ā�����e$S��I���m�%�#�,���C
���ki
I��x0Y�+��ڴ��P%�G���Ca�P���m�O����4bu�ΧZ��]Ƒ5��:H]���@��� [�W�t%;T�����?�����;&2�{z�'���p.,�	{6B6��)�'|�el'`�����	���ֳb�l��vÑ[�P����fc������*6j����)�\��L�u"�ݠ��������?�8z�����QhMe%���t'>��2�W�͎dc��D�|��v���R�]l�dmF30�%�b@<��?G����C��W�����6���ͺ�B���}o����ަC����~^b�v�6���oʜ{xCm 35�j��������=�<��C1/��[9�3J�)�k��4�ǣG~�W.�\H���k?�W����Ȟ��ᥑJ�p:�߶1��-:���$��cJ���:����U�<Z˵p��_Q$�縳��R���:�U�Q/��u>F��Vߦ�������Ӳ�T2r�Zg�~��� �5��M���T~f���J1[R�*5ć��GF�� �l?Ro1TR���ǸG>�����a�h)�m�r���l9���)�����E`l��mN��$���% �ǔ�i!��YP�95�li�Dy��ae���zk�%�'�����q��0V�m,
"�φki��&荚m����gExMS]2{yST�i�1"~Ӯh�\�,��R`�F���"���R�`�G)|�b��Vg`?*��ۍ��o���������˲.�!�� if)@���!��_L\�������i=��:Y�c�"����;y�1P-ߎD����ߚj���N����*-�T�kD�_(��0WVo��4�*��p}�ء�Ro�(k�J����2�D�r1/�L���N�\�2�!0ui���3m.�R!+Vͮ�I��ӏ��'`a"T�HT����i�'Pn��}���V{F�I���
]I�_�-�a���Ĝ�c�L02�Y�����K�(� տD�04藡�;��bj�#���;��2`��9��nd1�B5MZ;����5���D����t�v|��I��Kc�s��_j��d�#���1�vɅ$ 󵏳{4���ХM��m�Z�ɉ�-H�=N����c: ��������ǯ��l�4�2l/���ܳ�Lj�ui����:�a9n��]r���K�%�c�Y)��s���ߥ��NKsf���L��a���f�����)�Gsݿ�a�s��������[:%&�BW�0��x�teL6�L�&�;l�*�B�r�G'�\U�)¼�]��5�#�ܻ�$����2�/����3��BP���/`NB@��,]0W��=���4I�d���p0$T��%s�f�����
�BH][��Y�8�?�V< �T�D�!^� �_ڡ��s�l�z��c����HS*��S��X]
 �9ӟ��S���ẗB�Z��6���M��	B�����f�Htp��HC��B��$�����`y���������e��.�AC�= 9�g&�հ�X��-���A�>��@sU٥��v#i�j�8��^nK�ձH~B������v�OAG�'57��|����xA�#<��X���eM�]B񠩈§��^�{?	��N2��N,'��c�g��ҕ�2�h܆>A�W�}��W,�ߛ����g���w�`�?)����y�D�.�{'��4F��c�pKa��N-�*h�L�ׄ��z�_�!d�`1�!ʢgA^�L�z�+��~�
L��?����q��Zy��~��3V�hO�����(����h�H΄L|u�8�������9۬q�q�(2�jP%���ү�FPL_���d��*�Kټ402����m�73����ą[�hTTm�s�:x2��S�C��iw��.�E��9j�3�՟C��`mt>���"����R��C�jPE�Z/�C�G��a�s���zWw�u��α�O%�ǅ=�#���6r#�zɶ1gs��a�O�LA�����2�&�{��u�g2��)���:O=	j�ڳ���S��b�4ƃ�Mһ����*Õ~��oiLi�2��_h?U�k�uְY�ي�)Vq�S������i�����82<���vDr(3 ������4�?&��PX;I.�-nY�aB�!�oIq�/���U�"S�*}Ee1^��';�z>wt���ή�&�/w�L�^IG6P��Y����^�R�/Lz5��x�{W�L�������Fl�}�L���s���#�N:'���p���J�v���~��,ڄY�sK���ԁ�jN[�1o�2�E[�Յ֘��!$6�vq��G@�=p��ٹ��?~�V�n^��u���g�4�2�]L��Έ �-	����� 脋Z$pHDY���M+�&
φQ'P��ene�2Mt��7�x���E8��P��ܮ ������H���Yæ%��S%2�I���F�b����)d�2,�P��9&�s��K�E~�������C �Ώ���ԥ��x!��'�< W��<���X�Ṷlo���Q�	��,�cF*s�{Ӷ��ܒ(2�^���]�h'D@�ݧg�%p#�k���#�Pa�ם5~� w�%Ǿ`3����_��׫ġQ�SbR�}i�۔l�JVlX��3��#-�������:hb:���"uً��A>|�V~h�h�Q��2ҷs�����e\�le�&���߫w?�Ĩ� �ht����E�q����ݠ���-�~;P&s��ī�0�?�@IdWh?����f$ȿ�Ji��N�n×t�ԩh�>�&�E�������O��,��ǆ�I�����L:���Ĺ1KZ���m���@�O��^Z�S鮭_�6���
II���ڇB���>k�wT��I	M�vv'��(i�Ў7�49^��>[5}r�O����	�-�ܰ��@��̳��c1�R�u�8[����X�xI�kD+���5������Nw�wqx�;��~��{�����F���XF��⯾x���l�rǖ(��*U�����|G���sCi�m�(gF�%n���(XPR�Y�b�)����8��(�����!�0z�CGܯ�KΖ7Lc��,���fx� �{hA 'A�@3Q�}?�&�پ1���E��J��U�(q��������xv/�vI?~
��^.���	3L�p���lo8e!Ώu��/���((ԔU�K�y���� ͥ�5����!��E*o"��Z;�g�s턝O�9�	h-�$P��.��*���P�p�%�B",�qq�KE�
��⃅�$X��(���6ס�D`ZaB~����	ն{�]�K���#��C~�C�1Df��PAr˄	�����?�*�cʴ�Gc�Ǘ�ǩ6�T}�wI*/D4�#�P�8�j1ҷ���iVrܛ���%!YE��O��Z�z}(�~��f�P0�J�IY\�gC��n}L�������x:Zx�%�����GP�|h&=`M�wyh�o��r��4�qpP��o�\U;)*��k�dN�w/Ӓk�w}�5&k��_��
|0���6��hG6õ�}��.�d���2��O����N8z�x�zߌ�K�,3��GV1�lq|�:�<��|�}X����Kf��MY��>#
�.@��b���+Y�@;�T�;�4"D�46�z��������Ml�Ƈ��emr9�e�o�
J9�qe��H�i�/�m�\}�	Ս�ϯ�F�d&HKRl���Fp��IL{��?��� W˘���J`W����H8�Vbxl�I.,}V"��#�*-�"J�CIuyy��M}vc0&I�Nhi��>���r���z��5��|m��0j�g�ri�ߎg�GB:�z�?�y&��n�+���;חO�-S���H���j���z*��!�d"*�'(sr�4+���V;�ߟ~�Y�2�#7R�W�#���i���"�SSף���9�F��n_��?�� r3t�s#f
�L��V2��7l�����䆠�����o�P�ä8�E`]��@���)�L���|��F��ė�J**�e@9 ��}+����#�Y�)�6� `* J�%J��2EY�~O��Vx��}��B�ۋ�|v�A.�4u�4�=t��:��-���P��@ �UlLȇ��K#�����PXsX/�G��)�b��#��߲�)���l�����5�& ���Ф��N2���8�C�૆z2IE.u����IAlx�X��;���x�j�W�A��&�f�n�[�3 ������#���92т�>{�+W�%�������][s�{����x�l�^�����d�#{����琋
�?����[U��֞I;��c�}c��:�6��S��ݬ��B,R,�p��J���
�	��N�г��`�E���������}���G��3���\n�+s$�r�24l�D.�P��,��4(�z�2�?�w'������T1ϣ��%G|-_�ax��$�WZizL����ֆc@9'�T�'c��L��X;��#�0��s�[�\Y�%�P{~"@�;iΤ4��\E��dV����d9c	��c*�݌�Lǝ�E�)�vƥA���lK���6���[/�5�s����L��*?x�w1��1t����� ��)lmi~4UQ�������M�ה9Ʋ�"G���t&�R0�Q�z��� k�e�­���x4h��(T����@�%c�I�ܭ�:�G�r��Y��K�&�(�[��2q����ȫ��ӗ���e�$gQ���D���ȸ��������d�Pp�_�y:tQǪG۞z�x3g+�FA6KI���k�ܹ�������	G����@h�NWJ��7���e��D�vy��n�\P (A�6K�<A�Č�� �s����f�1��M����۔[�A��`��P��	0~�e��<�h^ZY� a�u@X3�$m'@��`�������SV%���QSi� ��q�!1�|��-y�:�����+�e9�T�^4�Q���Ut5Z:A&�y��`hs���ŀ7������#�hWB��G2������*��S�ʕ�W#7@�R�os�&�{�d$�A�@�f/e"��.�۾�8�����i{H g:���<����.�&�P�e"��=;y����)�3�7<�a*- �A�����.��C��T�N`�M�g��TA�8����(�o0J4ߨ����]���(3`)��|�DE	l��J:2/����x�v���;�2���#�/�d� ]�
��Of��}|'}��
<N�1E��o�M��4w�ոF���뙷T0�-{V��@h[t�^�7��m6��QQ�����X�LdFN��V��Qw��la�n����l��'�i`96�{x۬3_�Lg%]�B�K���e���`;�0��G�o(�UT�hf�z�Bla�;��hϢ���}�(�m�h�E.PcQ��|�:>� z���zC'W`��|]:6�w��g]�=u ��j�`�\-�ф*H1�~S�H��K�A��;���wZZ},Be���IUД����s���C�.F��5� ����"��ͱ���X(����\���n��Eڕz����M���㔲�ͧ4�5H��g��<}3�|?�]?#qg�#��2k�[�ja�x����^�jA�.�2]�=�wV^�)�H�#��ѭfm�#牠�b�-8}��D��;2%�	D^TQ�f��k�~�7�"��A�7c�V��e�J%��u�=�2��9^l>���:�2Hjw�R�|��-��`�9UΗ*'w��ޡ��`Ӻ�'�-�a^� �	��Gm�d^�����р��*�(�vB���r�f��ZCK���Q���2ʓ�_"���BBG?�-c����ͭ�J���z��#]DWX}���׳����/��z���	��ۭ��&wZX�ǒ�> �i/~C�}i|�V���;���������G�W4m���LQ�����'�R�A3n�j��K��H�A���b٨E ���@�o�\��w�yɗ[��}�.9C?���\{���S>��,}�%��y�Vu�#Y���=Ip�Z�֖��c��<���)�lȕ$87x�'��1����HC�151s��6��!�=IZ�I�E�]&�|��G�5C<�`,�M�6�l�_[D�I�ʩ=�Z�?��)��fk�~gQl6;�:��rV�%���2��A�gx{u K�ClRC[#J�]
�� Q���C\�����2���K���'#���+bjJ���to�V�!W��'��6�M=�X�Ҟ�e�
�I���C�h����8ZČ��{�X3<����φң�����=�j���D^��9X�^3P��כ����B(�L�/,Tf�7Π���aO�5�_C7�Z*@~b6�s1���$5�@"� ~�tZ��̠MM�����W��L�tA���]��̊<�w�Q*H�R���9f�2�ihh vd-�>��f�n�-d�������C�>��.`�kQJ�3C�[N�!`��E��ց>�c��(ȉχ5�;�V�1���y��^o�A�$����;�U���8R㐳_�JI=��`�x���[^P���.�b���̹�!�v�:�RA@i�^��Q��N*K���SjW�W�"u yT$�����H���׵`h%���݃����s�B�},�������2�(�c��T3nh8�>H��'�U�'8"0I��}��v�~%j�=����	�[gs���{����:o� �R�U��7(����䴓�[�$�k썤	��z{����)�(q9-��?���d���6Y�� !W7��}m����N��P�n7os�ݔ.Q'�9�R���uAuq�e`�]QK��ɱ�ݥ��0oo OS��Ac���А�9LD'�◙
�لH��&��_�7�xi���	��	�������T붷U-~T��x�@��Q9���C�<��!����ĝ��¾
9�
���dU�QͰ�|\Zӊ*�G5���~������D��|����q�طg�ɏ��dd'��9��Br��	FH���Տ��,�5�҂Q�+�j�6ř��L�~�_���Φ*`~Ww_��*L:_�����AF8�X ޾��{V���{e�ס��Ch�O��XƼkw���D�@���D� '��v���
6}kN�y7]�;\��$E��C���o%!F�ze!{�B��)E���������#˛� d�	�����I��ͮv0���s;��(ݙ��2��
p6YWڐ&�7n,�$?�\ϥ�ı� `�,�*��v�H���W��z&L��3E�f�U�,G���5;���ա!�#�s��L������K?����!/[��{��P1\�5��cP�����t��~����C�uhsFƕV�M��䎰�9���e�.q����e�b�`��g��I�&�]��$#�v�m��KL�����x��.�8Y��m�CV_n��p�3J_Q�[v�F×����Ȩ(��}�&�!i<&^���1�j~��hC?2����D��['`����(\�h���Pb�ڑ}f̐v���)�qfR�4���*��eo�k���Btg3jӻ.������n ��v�,C��W��ߪ�˘���� � yQ7�f �l����j��f>M��dY�����úi�����tT&Dʤ�Qu�|�1|�J~�%U�|(H'�?؇]���*���$�Q��>���&B��(j�90���g߫C����(��m�'&m.�H>uem����^p�g�x��-d�b��@YLQ{��N�N��Ku^2]������I�N�N8���*<yq���z�<��w���\�%��>�r.��Le���9l��yh��w�t���8��Os\`�y7�q�Σ���vX���EAί�4V�q���YW��[��7<�F�UzM*��K`P@bh�#��{w�F�B��?K@k���PMrV�L�	,��6j/�-�ъ��>�,��;���z-���w��U�x��B(�@��ë�ao�F���91dD q����SdD����H%����B-����!�%�Z����"vn���'B7���վP΍�r�0���w�vK��t������^$�42�G�@�?wɱp���Ģ'Q�[�ݯ�*�/b{��Gn\ ۼẪ8���q��n���ǣB�ߨ�QA���{�����o7����s) �4��<�^�6���;�5�b�<�Ƽ1I�U(/�A �Eآ�0;S�6{�t�Ps�A�$�]u'֤&���q��ZDL@iu�h
�������I҇���G}6CA!3��NS~�)�~�҈�J3?��
�/�,�k�0�<�D8�/�uKܦ�Wk�Amk5>A�I��8��B|#@Tc��כ�ڵdi��$��8J�\o��_�k�o�-	��j�SVXъ�~)�=�~<	\�K5���d���3P'��7r��r����P)��sa��Ln}�_Ͱ���~N$�8�M'�aIb��������B4p�i9�IK��v;�x��	���=�Y��8�
Gv�D�z�:�����"��%����׺ �������K:��ةAk!����E"J��\Db���̱t&��*����g�,u�MjG�k����-��8���T�Mkv���DI3��)���b,N��.s������ ���j�=s�_�����z=�~a}��m:�#9`��E!�O�M��2v	�vA���O��Re�n���.!s�X�<{�M�l�K�&*@����/�vd?=5�s���W�k�v�E	#���@�7�2{ �Kv�6��3waP�׭(����y��d��_���y��xō���=���u:PTW��Dj)�����ſ=8��Z��]������X�Q�!?~�;�ǖ�$�om��H�K2��@d.��d0�PJ����ę=F�?�=�W�'���hJ��K���*���1��o ���%w!E1��z�Kb#�t�`3�A)h�6_/���]��=E�vh wc�L���m$=#S� �*ee	#x�&9[E�Ki���{zD��.\����["]_C%ަ�J�tp�B���5������ �3V�����$�a`��\J�j2�k�����P7��z�d��=	M���)��[v�	x�I15pO3s�ũ�l�
1�mƱ<J���+�����o�E��ue��g�al�46�n��i��:� <��	TS4�ǣ�TI�^`C���ܸ6[S�-���	��sE��='i�U}��v�?À�#Y=eX�cm�����e�k�H4� ��w�	*���{ ���3���'�bp�������-d^�@ؗ�9=t�c�y��FW�.�Q����t"Ř��ơ7�%�����h\�����p������l�o���&�{y��Ҧ����a���9���RK��������N	��pg_�W����Oz���Y�̙75R��i|J�:P˅�<�c���@q����-���ׂ`���&ަ0����"3,5d�{0�A���Hmu��@`E�vewD����c��2ItOq���4駪��������Z���\���TV����Ds��xUAl��!�(��弊���o�� ��jg��ѴxU\��z��˥n��G}'��D,����d�fѫ+�h��%����0ވ�s�+��9�"֌﷗�D����%J=��n�f�=�g�^JS�Ԕ7w��j�O�zZ��S�a�&K�;��fny���7��f�6�����s%�傈�
W�sy�H�,M��E�Ѿ�!O!��P����.ѓu�lEeg��2=��&�Jq��ǩ� _k���F[,�t�)�ِ��OL���	�\爡�|Ss�>�ldվ�ElJ@�iؙWRQ��I�xD�P�"/���^�<�t���a+�yg�&eG���.�	����M@qu�T 號&�C��<��u�A�i�Xr�xqoP��
�c�-r�)ǜsphy�9I|^����ue������e�� t+�c줠��%�\)ξ���yD`�)t��i�v����w)��K�s�m:Xr���Sݻ�'Ӓ��p��Diz�]s�1�tCЋί�q=*4�N�[ٵ���Ӹ��N������=
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�ؚU�Uj��_� �~2
r��nA`|~�	���11G�)&�3�;3��zb�o�$�[���!�����3�P������LXk�$�=�uze,m��I`��
�`2�:|7��H7*���haH�x���6��z4��Ċ��PgO����჉u$,=ğ�m��:`�� m�X$ɭ�}�=%�TQc@���r����.�K���(�@��
wܶ'2�6/,Jւ��Ѥ���xKYN�g�;�2��.��5���(�l7��'�S~�M\n��t���(�Zõ���c	:�,@I�,j*�j����j
�Ue�D���"_�2��z��HMKw-u+=��
���P3fF�99�>��'G@��K��r3]����^�d�\fP�?��HG�t��M�f>F���T>�e6B <�A�n[���U��R�f�����y��t�
�V�.YR�5/�蓃zw���A����I��NI�ņ^�Im����!M@���a�����`{�S�u�Qc�N�7ǭ�Kl���k��7��+�(�A�P�J�o�#���?���Ix�vU�����{��E���c��\a���U���a�z�N�ڌo {P�>/C��)p���n�$���S4Y�?�>%T��)&/�1��-z�GA�S|>{ �Wiٱ'O�H�����m�>�k�E������v����^R[Qj�����/�
E``l�5��z_U��,��S6QQ���;M\Xp��n&�{��+����O0�\nv��������C��*�Ę)��m,�����/��;�c�ah�~%���R�k����	��	!�|��*���/0N{j�J���yU��p:�0n4���|���,��Mh&{O�L�������|b���F{ ����Xv/<b��#7�d��Ȏ�>/��zn��Ӣ2)bA�Y�������8��&���U�^HOe v
[�_�\�g�S.D�A���3�%=�X��q��}KAZ<��Y���{"�{|�P�C ���ȇ.���MI�Z1I���FV��J3�0���?�pzb(��u@хB�hB�q���0�� :��1��$���pّ�D�UL�H�"k{�Usf}(L���#]�`��e�(7�0zhO�?Ƒ9�`��9��^LɳzQۡXo�[��j�-/��X�qe�~yRw��ʚ��/�U�K�^x��auv���8�l۽]4 Y���O��҂����*H��2�$��H�=��5����m���7�a�ZN�4>܆<Z�9��U::FU�SYr){> �mWS>�iG[W�P��-�� �c��\Fܣ
jm�K˞-Xq@�k+�1����LX���Q�Ѣ�i��g��V��zE�Y�X���y�p�\e�I��s#�7}�����J���ްum-�<$�,̗P'"�ٸ���I�=S��($b�����-���p�v7bw1$�78���naΫ;�%&��I���&��5�F!��OD�N̓L0�
mY��|�T�U�v��f8��P��w�I���Q���m�_��֨Ϙ� V-��z�1��s����t����w�T�lp4�{LLQ�����v�V�J7���>�I R�N�w�����2RE�m�C�t���S��aæ��8���R�
L&�\O���`����w�1vl�p�f[<:[�ƜX�8�v���Cy�-_b���K��U����'�9[g^,����q�KIq�=ζ�lF�3�����Ә�w^#[��O�1�F�l2���Eh'T�N�����^R&�5w�J����si������#2���Cl��ː�o���C�e�oRM:��؎����*�ί�0͆����W n��7X�o�����灯��G�A�^��+�Jx���k#=C�A�6�J�5��VIg��BZ��h�E��u+Fw�;W�<�
l���-�<�L���2p��3m���zUy��A`�&��JS���U?�\���`[��D���mE#��>q��ۑ9�lG�Qb���UD
,&�Ċ�����Rv��H��ZެZL�t0�z��Mj��Ck�"N���Ç�/��ᕯ�K8w�����/|Oj�]�WM���͈^�JL&�	�g�{�c���_�Xt�o�g̙�_��W�f������P����*c9���![lE�"ޛ�ѫ:�f\� >U+p��ɰ��)���^ט���U��4{-�x�7�wY0�hT�����p���0�#�&v���nd;������b���g���N0�,�>n���at�"�t�k�x@�Ly���*>��m��%�6�0�D9��6ʄ�ZW���t�]dbA�(�3���?J�~g��D���|�u{�&c�����'�A����ʳN#"�0CK�7����%c�Ȃ���ty�q��[�W���K?�t�ڹ��BG�Dy�Qv='D��%�9}���;�G�"��ˌ�v����h�'R���ƃu �I��@��ڋ�&Nc�࿹a������񒁔N<���� �`�o>}b׀R8Y�\,�ǵ�2���]�)��!����@����NVo(��9F.1��|���)����4����ڎ��z"ܧم�,KC<�u��c�
r�w�L��Z�w�����TS�juJES:L��� R*�(&�א/�קn�zG&m�B:/�e��������`:D�w�:�F�J����^�|0~��xu����C�^��:��8rە�y{k)�i�����NT�<��Bl�F\~�"��<h��qv�e��F����/b�:�d��|m�G��>�O_vp�5:{��$%{��YƩ+��(;���'x[Iﰥ� Z__�=��� �ǘf��0�0���S��6S��FA@�W;��J��2��V�6�����7{z�
O�����:�����ry{.m�o.{O�Ym�����8��5������-;�C�M�B������o�� �ř_�����T/:2�Z��k��(UAp��j�,�@�|w��m�)���gҪH3dP���6�e��cgI��k'���Kg�\6eLU�V�k^ylg��[��jh����Q @h��q�'e�ȡ���V1�I��*�xh��o�c�C4�n�h:g���H�DJ���M>��i��g��}�2�Dg�`�P��6��o�!VP�_���j�39��~Y�Am���aqWX�f�l��X�����W��ɅoAK�a�ק�D���<��]3���x�\o��U�Xx�u��;��_����c�J�6
q��V���7lvD����NR�4hJ��Y�J���!x�~���F��`�R�R�v8NE2a�d��<�ȵT�.a�A\4����JIv�ij�b�� �3�K�'���&%�O�܃�@�B��:g�9��9�����Yp���\�+��_'�i˖�	U'*T]9:
����/^�
����6eA�P�~�YH0�����0z�]x05���Z��w� CY[��`0�']�f���� [[���etN_ 4N��sP�3��9^��6T�׊J9��� ���k n�5 Y��(M>�usf����k��	t�����u4�{��>�9m+��ڥ��B��/�9�)����q�[H�DV5�|��U�N{~1�U��.Rl#D�� �بB ڸG��VJ0�|c�1\�@���4&�����0j��ł��d㿋�zh� eR���<��G�0���c�����it&D�,K0)�� z��?q�G8F�^��3��*\��=�z\]g���������94�c�JɃ�T�Po� �%�[��&�#Ҟ�ǋԚ�|�o��Ǳ�I]o�ɢ}��Y_z��Xw^�s'^V�D(�_2�M���";G���' O�Q����Es(]�t(ޟ}�i��TΓ�����g����cJ4X�Lڏ�ܸ�]z#,V�<�6�V&A���lx���;k2��H��	ޚ�k 4�� �[��u�Y�c�2���l���w�m�Pc�cO��m�
�%T��$��",��\�^�&��GY[��Qmf��U�t�>��P���66�|���1�e�T.q�Y�a�f��xx<�6\�˼�[�����.�1y׶�@I�PMn�f�CKo�|��mӁY����V��⭝ac1�y+��`\%���i�?��#B?c�������V�8�a� �ѝ?p/ ��PY��1�`}���� �z��k�^�u��$���oo0[��6/�?K�H@����[~��qu=�^{d��q+��ҭ@נ]~[
�^]e2W�w���Q�٩�I��W@�x��*X�A�6�;t����j���;&�,��-�*��P����D&�(�H��"l�F y3�,�F4�>B�������`h�˜����ȕ�ߌQ�τ0�|���w��o|�_���Rq�"���m�C���d0�[;CMF�:1CO�&�Yp�=T�r����z��V�-��`�jg�~�9��cw2�sU�lxTAbM4B�j� }�S���i�'V��հ�M=��ԝۓ�rD�Y� P�*�ѝe�����R��U�dz�+�~������pI��g�B�H!��<�zŻ}�.�su����,����sd24
�Q�0,��9M���z�>�kMd:>��K�挤f�b�T��H�Q�l����m6�N�Eq)�r�N��o�yF�*�O�p��pi�2Pb�͘O�&b��f�������A�{�2�ĊK��4Y��G|���#2�LG�n�qM}��渪OMfmB{q�A^L�r��!Dz�#���-8���T��C�L�І	�#P�d������s���)�I���T	̦'���?Í��J�m���U*�DS�;��f��v�U��Ķn��׏E�������XE~��b��.�T��t�)�Og��9���g�#+;߆s�r��=4����msw�F���d����9rX�y���Wʬ�s&���T)Tћ����:�:��,��	ky�x��Og�J��{�дܗ��L�H}��/��XY�@��Ʊ���D�v��ri�o?��: ��#�!9h{r5��`eM6.֊��������.���M}����xH:�ux�C�D>)6	+��۞F����_���?bH��S���d�ї됞��c�����:�  jj~u�Z��p:c���G1+j���H�:#�q��R�dǋ�n:xQ�Y��5�ࣶ��]�(�F<O�d��sa9:���/H�M@�!⊴+��Y�評��sǔ��h�}I���WƄ-۝C�w�.�
��� ~���e���B�{�_jַ!���x<�!�7�Ľ�_X?ݬ8�8�ϼ/6�7���F(�XlMe��@���L�[M��������� 	D\��g}9.��F����W?V�.���8�2�z��ɧ�՗���D�7�C���H������I:�����DbP��מY�=��>����Ti?��~`h�r�Y��	W���B ���;�O�aY�'ʫ�����R�¥��p�Yv�ďzYڴ[ ŷ	�5�O5b�3������1�|�(En�S��kҎ �j�/����̢�d�G��O���i<aaK�x���)���w�IYQ�1#F�D[�^5&���:�76GrY�bzm�J�cV/n�7�s7����6>�w\�a��S���}p������vh�{bNJ��B$n�*��p�|yx�=�NL�͛����,$�a�(}�	i$���ݐ)�⟜�Y���XӍ00m�l�Fۉ?�u����j �� �0�_�B~H�K���?�㒿U�M��{��*J�0GC���S`�]?@�h1��-��ܢEr6VĿ���c��\�K-?Th4�����l���o�Uc�r������Τ��$?�WY�xŇ5�@^"	g�?�'0f۟PA�z�Gh�5����9K'|�7�����-���O���9�D�H�r��IJ��p%�;�>��3/�"�ޅ�ȏ����9����wQ"~O���/9�� ��hF:&g6}�Yw:iFG�*�K�0��mS'آY<�p_�κ��:��ב�C�P�,�2B�����xz������"�͋����#��4	�@�:��3������G���4Bv��tL$+�h�޸2��aQ,8�9bs
���cZ>��
C������"d�A?D�Mh��j�֕��SY���C�9W�$t����Oqړ�Ž�\��m��:�{!�Y�TzI4�b��!��ld�&Z`��-�}'*|�F\�FK���2�5_.9Fz��"�S�jNߥJ�
����ł�k����y�7su��pj���5�nf�j|Thu�Py������x�O��ڊk��@
�÷�)�ğ���=���A�2�w���#t�����d��y���D�M ��x|&&p����xi������>��Z��U8�n��*R���%�gkc�H��8;����J�ֳ\�>�B��Ŕ*V?����D� SY��~y}��:�~��B��yl��5�Y��O���&� �(�7�*�m����@�ҁU��j���>;VG�I�	A�נ���7�x��4��xte|ypV��%�cu�<�7�y�����k��p��
<nS�7ٮ%ş�l�m�����\a	���m�GaХ����k�|�R�|՟A��cJ�:�x?�kC�΁�����ҳ����첬?�Ͻ��b�u���3ݶ��m�2� S�F�q˧�Z�ժ�_{ ��q8��G��no�s��5���;�	�_��^xݽ�{2����Y�vP���M�^$�2��h���4�z����5 ��X�JM���'Vv�׋j��LP�1�V��AYO9o3��A���aZ���!^R����>n�k�Z��Jp�-����Aٍ��s�*�B':�^�
�����0�� I���x3�����3�e^e�xl��h�!�
�w�m&{����u2�XO� 
��#'��V��"�.<�E(c�DH���g��wĜ`�:H��3������y�дV�m��O��!�����_B�ye�XD�(��:ʨ!cL�N7�(&�T�)��:h�o����ҵ��MB{市���b�}86��>��#��t�ұ����<n����&�:���L����o�+s��̙o.��,7���Vm���b�~����[Xi�xQ�l�-~Hh�TU؞r�yӉ:�����0�̤�!4�k_���$��sr���땢T���*��&�{��d��7�Cs#��H�l����B�S�!x]���ͱ���#%&i�

�h-5g��e�$�U8�)=��:� �Ɍs�`pI\s☨"l.��6@�f�&��K�щ��>j�F�,蟗���kz2�E�V��k=L��c�˃%Ս:�]�8��f��Y��_*[�6[�j}zu�����Q;[B���а6c��;�#�+A9����"	Y��^F�)��F�O��!u���d���-1���#�U�_�Y0�����X����ς���P��R�e��<��-ٷ�����pR���Ve��N&�3�#��Y���fJ���F�����fu��Ժ$5���惨_
Ɋ�K��J�ȋ��� ݏ�vҐ�a5(t�%�a�;����9�[)��L�e�O0L=��]��lLD�dH_���s�j�Ls��j��	�kJPN��םBa15`��ܶu[�z��橬�8��F+�
��^��"��B���c8g�"g�{Y	i�a��{��%�f��.��N�LN?�#�
���J��N >�2�p�=(��=C��=��|��rT��/��~t4�<Ċ�x�O�˺4l�%������95a˷�����sp��NR��N�wG������J:A	�SE���2����4�(�1�\��g�YRІ��Q�+֢�ݎk��+@0���s�-�Y52!��7�)`�ы�H;�i���e�A�|�%�F��p\��1 ����ǌFiP�2�V�V��=3��9y��R�ds�9۪�EÀ�V�B��/B�t�?���¸�~�!��K`��|�#���3Ns�0���Ayd��wL���{���'���Ri*�S�cs���P���j�?��m�F6��yw
N��:�TTԺHc��⃷�YO���:�ޓ`^�#Xg��6O/Q�Z�m<�wL�;7��jT�g��Y��.}ۢ	�ȨA���EGe{w�݆��#�28�Ҳ>�{W��My�d���gQܮ�������u����)�4�ʎzb�Q�n3�Q��q��6~QX?@�.V��W��i�2IK �*ސ�İX����G�jUh�ҺE;�����V���L�	!����::����eo�@��� f������1o٦��Rc��=1���_�ԍ��ֿ�{z Q�H{fB7+gחևw��	G?ݗ��R ��Wݑ�zW�:���ܷ�r	+�^���kM�c(���!�볌/�R}`~[�l(��dn����(i]��Z��:�@�T�pR��J�{�b(�Q���Y֖�Q�>����T�Q�z6�I�)<�$iG8ٽ	�V�$���ynF=G��&��G�Q��u�IQ�b7�}��!�g9����f<r�O�ՔQ���j�����1,�-�)������t8�%�t�4�+��u��GH�6�|�5e�]�7��7����)7;�ѹ�t(!�R��<rqfl�q_�n�Bn;E��9��mk��1U+����>�Mt���j�䉮�-|Y���hhz���-���u"O�o?����rB���/4���F�~~k��T1��a�65��H�U�Ҋ{�V�0_Ui)��:���l{�
s?pzyO7H*��3��Y݅�9)m?J�哓�[�(��iT
���s��7�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@����D�A=O�"��.i
��f_���Z���B=��Pe`�b�yi��I�!��Z�)?�!�4��p������MO���f�r?1yf�tQ���-|��3�5���n*��
T���Ϊ�a�����r�8��A ���2@²<ִ �z�KO#jD��]:=GS ����Q�Ƞ����$g�>3���|���P�8�j��`ob�m\�DM�
xrHq��:W�m��y�k�U�� �-�|��%!H�K����,5ǡ���N�
l�I� \���̷�9���.�!�}�f%6x��%.,��E_O��P�gy���&.��|�;޴{ᨧ;��xx(��M�����e�_�w2(A����_{_;�˳u)M7�x9`s��qE�=��� ���JSy�0?&$��Y�������@X��`��'8�cGHJ Q����\u(3��P�<�kd�Z�سU�Za ��(m'q�NN�~��u���r�嚴�@����14�uosc_���!�I�_3����=#�MF~��u���1eLvBf�b
��t��η�d��Qփ��fHt[�-җ��Ϧm.~�)����u�=iM��+C������ҧُ�D��PA:b����6������ϓt��ez���la�RF֗��:I!���Q�P.��ҟ�h�	$S�5�+GZA�n�[�zWu�,^?쑶D�!�J�X�8ɑ���g�T�%g��3���-�k	'�%OMd�9����&����k^�� _$~H���eZ�©��b��Ќ46�m�L� ���BxA���t����Li�G��ZZ���amΚ�����%���s9w�B1FfN0����r�;��쭧�	��X�0'wVPy�{�>������&溵k��)"[I�ԕ�Y�Oѧ�$�2i�H�D�
s��&%�q�^���\5@T�3�����tjX���A�-������)��]�W��C^�wl���D�s�W�RT��|�P��✕��yyvc��ҭ5m�+�u�9�>�ZRч��|!B�忝q�:��iH4���k�`R�_Ό�d�?^Ϸ4dx�i�%p���Z��h�:��άNB6�|i�͙�n��rkۗpdH'ж�¤����+��C	5aѶrp��T�DH]�D$N��Ek�r|~g*'N�8�����x?���%�����43r�����/#6�����"�qSt���$H���&��X��z�t߯�Q6` If�'� .�`)���P��V=i�^Cךł]U����*$�D�x�D=�k�P������q�'�U1�Qq�|JvwC�f5��輻	�f��Z��αڭՁd�]����R�����5/8�Mn�i�A������;x����~��0
�K���T�Xl��L�B_� i�ԯ�T&Y�b��a��%n6x �������~��8�>�>DD��	>����zj~d��'+��������.�����Ǹޏ��/�!��;ş���Ac���a]�X���4�oĠ/~�"�}[<����uV$��)ع�u�%&e/H&K��ʅCڜ�r�u��8�xDw��EW�`���hI3���2U��RoQ��	��*�����S�"3��m�.��8̙R9�#�j�/v����i~eR\wQ��JM8㵉�YE�k���W�q�/�U�W��3�ε�{,]RVӰ�8UH�3,��YH���[�f������>���J��n�\�� ����� �P�_f��ùز������)�?�;��rcܒb��4�2��1�:�vt/�6�ˆ�o�
�����T7� ,�ݫ��h.�`��f�(��>E��xh�\��CN��	�s���ţ�Z����I��E�7�K���vʖ���|R �vS�F� ��=2;��J��/�(�ֻ�4'�Yj�U	�YP��g�#[�7	�d�T�w�y(-<>���߲���>���������9GTw ~���;F �}�/��J�*1v6�I�ɷF1~K|1��5����(s���)�~����T�I�a��'���σXj�Fk��ƥ�}ʝ�|T"������M������J�0@-<�:tR��Չ �����\ǝڴc�1��WWyÖ�����H�Ct]����E@_t�Ll{�)wQ@>ؚK��i47�I��E�/A ]�6������L+�:�b�%VwiEE
J�'�����o&VU� 
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�N��ն�2#�&Đ��xm��D�[�=���Tvv����g�5���lphl�(���AQ
=���ٱ~?�A�1>��^P�OLK�7���8i#h}�y
7�2���c�UNn���:t�kv���3���x�@��[�nL�v�Q���<���Dxv[Gt��I����c_ypO��gE��*R&5��y�0�8l�6�hβ�r(�aI >��>������P���S�(�=]%��튇R�����/v	�Fc��"͐U��c>p��d���x�-��R��k�p� �LF��<�m@��q�����Ôֶ��F�m �Aƻz�j�q K6)�ŋP�������Jy��c�V�$��x����)���o88.�nz\��1�����&'r������������]&�����kf��{5琲��Dq������o�x��t��P��>̈́�-����!������l�0\����h[yK���M%���Q)���1lz��Q���6�
�@�M�(��䆅�`�.	pF��FeW�0ZaY��͊�P�dsK̯ ���@��}n�C���{�hR�hs�h�����$<U��L�!z�y@"ծ8�����@%��VK-!����DmCJX�gNOn�CUbTrjD����)LYi�T�EZ�/�L:�o�Ä�@�WG�o3��%gX�Q�g���6E�T0��
�{����{����!hq�� 	 ��t���J��ؼ��!'�ʮ��6K��X�a��Ec�������q�.z�
Z�^nl�;=�e��W���*7j����W�z��P�e~.ã`����k<��J����$�/�!T���-�RU3����+��Q�]40���/�8ƴc'<�?���o�T)٠�����\��������"��Ûq�/q�ES|r�ij^�ޞ�:yY7q ܋b�����<�����Бp��=�^���c?=�,
'] �.�����Μ:�u�'%kS8RR����1��݋���Xy�dp��a?d����L{$ӱ3y��@�J	:�Zt����O�|�*��fO6�Jw�l��P��8�C���0�,6;J�&-���:`���ݏ���Q�͉Gj��I�
�AEVVWi�u�΄gpV�E �F :CD�q�Q�,(�Cp�D�����sT�@T��V���J�w}+����#�O�vk�]�Ch��_�4�~�N�(�8��*���źxh�����e���;��D�HJ,���<41gu� z�5-?۔��#���'��{{����z_���7��-H�I�Zk��ɘ�+H���9�A�{�k�f�r�ߥ�����»�-9	]3�Ť9%����o�\�m�7���	�_����z���k[�*61?o�ƈ�Z.qe�.��қ50�*b-H��>K��7�����p�K��J)F����y	��'�wы�O�dy���	O�O�l(��㗮�J���n�,Ţa#�*A�J��p<{�� ��ߏ�����q0oes��w�"��޿�4�j�����(82�DZ�.��T���R���4�B{l3��RosΛ����V�]X���<:�ž�z�#��h"i3�&H�6��г'��rqm�y1��dy�
.h�s�/�K���~�=�MU����G�0�; ���Q��R�NG���W�W���L��5���suLŴRN��;A�z%���F$t�i��f�ͯ͵p���} �P���|��:��,j�ܣ����O�r�����&EM}XM�����9�ЮT� 
�{�%�-3?⃔���w(�o�12vԥ��n�c�MJć��Y��Q��wd��'5�-�0��_��,D`J�Ij[e�µ��A_|A��N�
Q�k�;P�����%�Yk4@��U����ϓ�dQF�ʊ�~w�|I(&S���\��b}���?���T��Oط�)�џ��;��|e�#�ExۚLC0���֞�(�C�M�n]S!/��O��w�r�K�V"��`wg����H۽�b
}��;�'Y(�m:��Tpt&;�4�+��o]`ڧ��d>�R��а5	v��y�y[�ޙ㛠&(1)�P�t��ơ�GWj�!/+�Y{���E��T��Hh�b#>3��Kz>O�A���|��=Мh�3�\�r{�{}q1O�_օ�,�㷥fM��ÿ�Nf�ѡ���dR����.�Z���������־�b2������0�3�\���L�u�>�K�~)b�%��^�>uG�)���WO��ŬȬZ����K?D��93�ҦTJ �1�Μ�'ڿk�?����nAs6�h�!�r��h�}���K|�A".m����� ���i�~0$Ur��(<�~VkI	�_�z�N�EF$�i7�E!��QvC��w��ڰ��>�~߆�Aʦ0̖@9���C�p�d9S������u%���i��7�Vn.!��M�C bE�K5P˃���Z�ԍ�X�M!�����0!p�]�_,1/~Ǜn�aֽ"��K�i�+�c_�("x�I��RS��]z_1��nĖ��y�#�3�ohq�]�	v���3�0v����|��p.��b�-��za��yk�B��Psff2��8�/F����H�{�{	�=�����D�`�Osw��`�'�r�v_���	����D6=D��m�� `&�|?��w9l��g�c[�h�Ǫ�e�F��õ�0E�͙�9�Q�f%D3˓�?�ڳ�pS��q[V��TP���3^��|�h�U�5{�P��&�BM-ZV{}��G�b�P���8{@vZ��К��K�����F�OfT����u h��R;�Q(?ʂ��zL��^V����J,��:��L�=�ce{i��<��z�o�/|p���3c�Rp�5[[��9�!Յ��}�9�p�9 ����L�T㗞�E���o aZ���x���n�v��<�%dT� 9ek$
j��5&���	��Be;�5��>�@9�݋>Ƣ��~����td�/��M��9�J�l<�1�G�th�o��6�|�9�\FW�V�Ǥ����os��p���W�Px1lTwvvdP�^�^�(�����l����������*'�DM��ȸ���Р�as���=*��ޱXY�-(�2��Q|���	�\kq"=�a{+B���!�����$�s��U(E�V5c�V�g�U�H~�{��t/����TK*1|�SiG<W�%(o��/ �F�E�d�g��FCO����c�7B�	l�R�!?	?��搬I��ot�A���?6ɝ�kߜDu��Q���7��fͬ�SjR!C>��ī��~2 �N9��wި!�Pj�[��Gc ��6��J�i�g��/��&��R�cTE{ۖ(H�1�����y���v�%<j�x �]K#�����;K$�"��h�@"M�q/�l�t���N������T�
��Qu 3��[�g+�ҜT_o&�?���.�ݦ���9��˛�3J�̈́:�q�?*q��g�@���7��?�wx� ��l�m*�( $�^a�Ό7o �������f�N���J'q�b�z%0<�)6cumz��j�Aފn,
�Id7tcY��:��nv���'���2�\�<���H:�ֿt���A%�;�W��]�/>��3�D#�%�@����0+�{�@(f�|k�h�bæ^��R�B��#O�l���U۷h&�[F��vP�@��h����0\�AF�-����.t���-����!2k�ܤ���+z����<��F�r9ufk�|�&d4����_���?��z����BN��/��ީL��g	���c�xC9�� ������Ԩ��lLc�r�Y.7�i�c�P5
��=>��tW����c��u���T���)ͻh�@5��A��:ؑA��!�Hb�W�lak�沙���p���;:�cWc����;@��a�ec)����u�^;-"t0s�j�}Y8�*�@T�!�/_��uRh�E�Y�����{�@���T.�ڸ�Mt�yvM�>k��?��R3U�O��Xl�ʙ��W���#G���M2&$ɴX��Sڗ��#���	�J��y�T�lL�)u*��{���<�c��o�"���ղ��pXd�TrH�<�5�FNq�/�� �L?�)�6�0 � W�OUU����t2O��@�ZA�[��Ex����MK
G:��]�L�s�V)���X.ʄj�\>�޸�EDbн�B��#	�i�4G�`��]
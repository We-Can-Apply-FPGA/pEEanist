��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i��������쀞L̓"�oܜf�~�5@�g4�5�	�
����,aeH>)�3+,���KԾ�D�X��x���ark��!��H�ҫC��\���!Q{���,�1�Y{�fd�wGP�n-���"����R�j��{��Ҏ쬟�b�Vji��a�a�n��젭Y�?T�K�1����MY�`�4)���Rg�O�C�p���5��la�Dv��F�EC"���L6�ܟo����{H����u{١l�hLk�輎A��m*����x�SN�8�F�S3�k�Q�͟碬��� �� 4L��
T���#YEQDWP\�9�ڛ��ܚV`]������dj��p�ETZ@บ���9�fފ��[�8�o��esO�/�nIӬH�޽�B�\������쥜��}ЕV�(5ø�>�����9��̮;}֎��R��C����5��Z�Ӓ�c�U���%1->�de�� ���n���Y �|/Ml'�q���d�l�B,1��˔C�B���s���`�g�\O͛a.�ko�]a�lY<w{x+п�q�ufg������d��-We���jux���Z��$fU��W:�%ӨOOcS؀r�
�Y����Ӿ;
�(G��/4��ХR9��y��$���G蜃j���4Qp�6��#���Y��%چOW���[��~�7�wf���R�4�4�rz��~"ٜ0���*��*Wc9�$������j=f,-u�����k��u-�I���6wZ�^����G���d�)]
���yX ��:��9tC)���r�|���!Řչ[2�J��!7�%=�����mv� �6�/�����D��<e-�%-�Dcs��i��A4rj�� rW���|��TB�EՏa���%��؁�9
$X0�_�1I/���d;�e���["�y��l&�.�� �t������rA���C�
�FT��$�*�d�w������I��.�=�����V���װ:�B�Y����\�o[?���r⬑gO���5���^W�T�C^��7��c��a�V��Y�]9��Q�ɷ�	���E�9KE��n	0\������*?6�;�(�cl��[kS����{���{ ^Q(9�\�����X�"���[�d'��(i���b1{��:oN�6�5��x��<ha�.s"�����}E�hqX-��hn��O�=�����iUo?�#������;�U�:_��;����s������2:�8h�I��y�b�)[ �t����E�˵��\2L��i�MHnFL�N��_��ɪ�CP���8��w�l	Ŧ��Z0�>SX��_���2���b$��!�݅��?�B�i�l	���������33Wh��Do�T��6<m�v~p�c�-���=81b������o^Ėͱ�D�NTw^`�<3�X�O��}{t�9$O�)���};�v9���)�=��δ�M������-�j��Y�N�P$��8�Y��VP����F��U�/�'T�������k}��wգ?"7F�pͺ�&�XЧ��΋z��EzRA&�ϷB�+����F��c�޷wa'օ��Z�p�A^�������~O$qi��qF�O�ųzG�HjIAN���;��������=멗���s�����{������6_v��2��Վz��ϔ�J����g3��u62O<����{P�T���U*WQ����g�%��cͅ�SU��vq�a���Q�\���1�2�M�f��j��e@ݡ�A'��=�fnd�������s�dW�ؓ���Jۀ����q�+�7RK���]�/�x���j��6nnܗ �2��+H����`��������5��@��\3�<�xߔ�f�^�X\g/����f�ɄW�m96�Z�wɧn�K�h'Ժ����}v�&�zT�>mxV5���~Ev�G�suD�r��0(�5C	��&1��
�Z{̆h�����<�(A�zE�P����-`l�>���S�U�m?7B��J�3ց�������P�.��˾��6�V�!�u�p���_S��XI�0 _a�gU	{歒�$̍Ԇ;T0⤻kr,m�1o��!h6;�YV�77�*uUr����C���G�p-l6R�S:5"��,�ĮI�!F��T.����n����V=�N�3�W3��^*5��=]~V�3�5=fn�Ȭсv�'ϟiEŋ��i�oK��@Л�M#))���/	]vZJ|����7KU)\���t��a#���}���c�-����kX��w�|��*�,��6Cd�"j]K��uͮ0B�&yY��\j�
���iZEZ���G�_����g�a�d���XV���X5��E�s��Y%L�+ئ5��D�=��
6��+�v��I톳>]���B��9�,�u���bo52��:d4�V��^��2���Յ�����yKo* fv���:F]H�T�W�_���LA����42 ��3�X��
�c�����%��8I��7�i� zt��.�ſ���9�/0K�J3���Z���:�PE(�8����5;{w����O��Q�Y?Cf�2����}*Ԟ��`�Ī��j<��������taۊ%�k�ŋ;�N�m�"����y�<��@��	r���Qz��8�U}�Ԉ��L�[Pj��;�ԓ�s���}��W7r,M6��
�~@��Ǟ�R�+$�\�T2A��� ?�Dk�'*m1JX[ұDPDc嶻��i���<Ў�M�MFtN+P�r����yc�����t;~fr�c��S#�TW���*���ڦ�ٳc�M(L/	�-���?�s������:��$�ζ�]����v��M+}~ٹT[�ѫ����@���YXϼr�ɔ{ 2!�D�f�`���q�΋G�д�8�*mҟ�4�q���3.
�\@�W���(�cq`J�Oȫ��.��/R����Q��s)ͳ�w��������gX�R+��RV�6r�EI���s��R���8c���=*�Y$�fո���#���$V��dUq���W���BnGd��*��p����h��h%���ލ�|7 ����(Գ
nx�c�������o��B��&�pOhۇCgoY-��T R+B�����?@xÿ�$#�ĀIB٭F�/ƻ�s�8(ը%2��E����C^����NY
)k4��zi�j����@�T���:t�y�]Y���>t�_H��?�찖1̷�!*���ۏ�߀^=\�s�����
0'�=�1�N���;����}Lw�(�T8�i��B���#������7�:�C~P��4�c�cZ��X��u�`P�JN�M�_�c
pe�9o7�m��.f�Y�\{�%o0Mrl)�����;o��~�>;}�E�	҄?�M-�(��[}E)E|{w`�r6�p���(�np����eJ��.����ne���&hK
#��	����ώC\8b�"l`Rf؎��;䁳�9��E.2�����i���N^����؎�gHg��=X�o9��l���T�乖����f�8�GB� y�A���J��������������>���r��#�.���)�DNާ|#��#����'.)�!5@��8y�"�!�|xfKL0���3��[z�εt4N=О)�!�*'��~	�Z��C��&��~��.2�{ ��s|��^�sk+K���%��5$�0�Q����D��n0R����o��D���_��"���,.�D�;|A�6!�ǐx{�d��U���IS������f��s�J�Z.,$�P���gp��ԁ��(P�@�M~�t���+³��.�2σٗH����~R�I���Q�F���e�
�#s�U)��T�\��֣� �ɧ����f�+�3xf|��*^���RH�@r�~R~�t�SMv;�Q��
"㝠��%�ù"/��I�[0��ϒO7�ԭ� ?E���_C:��|�+��lh�eU{v��=����Tz`(}؎�4P�9R�i[*UV�ı�E�}5�ըK;��5�D˥$��̤�2�v�c�<"6����MO�t$E�@Ϯ��<)���Wed��u��d�*�nC�= :���1��ya)�C�)�$u\KaȤifKy�~��d;�\j9���t�
.ǽe���sO�4g4�T�〕��m�1��s �:H���ǈ1{6]�Dk�+a��[�\oYD%�m����f���Z̷���9GrQ��F�,�������~���~y�/�s`dh�%���ϵ{���d����|����3��%T�&��`�p_��=ף�Ёc�L}���s���w>�s�i���nR͊�v5��|��K�2,��,��Α$پ����9\]�Յ��Qo�7�M Y}�D{RDQ>�WI��^S-�]�����7������ZA-<$d���ފ����~!��{�O�G82+I�>�.�+��a��O!||F�,�@r;��-��
� z��G��[�)��$�n��w�Y2��������2�'+��ܽS�,�S��o�Ͻ�}6�B���祤�;�r3R�A�Nы����aW�����u4�T���n�'m�{k�$e��)�
X[����2���p詮��I�_��q�-��|g�\�+���R��lУ�M�DN�Ra�^�_0ʕo�ٚ��RaS�د����*�%Wl)P����h�J�L�Q���R�zݙ��'����O{w1�\H�-i�U-L��dlmt�L8�X0n�*)��)�Of�s� W>+z�_�ےo9���I�j���^|��x��y�1X�~y��Ff�G"hme[(Ѻ������� ��0���Qn�(&p�V�Y�����f��D$|�y"��;g�&~dZ�����H{�(�J���pQ��TC�)�K9��y�u��Y�Lp����is���7��8ݑ1���%��_Kw>y�>��q{�]��:�o*��Z�<����<����1�<΢ [89��b�Z���L�'��V���N -����c@���H�I�.�p���N�+�10k����I��(k��u���.��"����F���<����	�ge���N�2ІK��!.��P_t�
ԙ��8�l�c���S�P�9������p��&���!p��?�E�cK�X���Z�E=�[^֞\��@'��h�������"?`^a�/.
{��H��2�6^��|�2~�2�����m򈫖��}�x���Y�H�b�2��v^^b����8&r?��C햺��󲗜���0>�bOvo^ə��)�+S�>1m>(����|�!kw%�R�%]j�!pg��G�-2���lM��@�JJ���~�����n���=�ΒG�(0�|���;�ీq�ԣո�^�h���z�g��)Co��D�="��r6�n�/!-�괊�C���@�u(�tVdt�k�-�8��S-͎ɥۛ����gu��tZW�A��Kb�Ϥ=� N|XdG��0QV-R��O�F?��;N�C�s��3l	�L?Q,�6s<w��:��A��i �f�$Q���B�.@,���ۧ`��%<(�D��e��+Q����j�f_S��}9O������(#*��Bbo�`K��v�y�jz����R��|h��0<�t��g�����3�Yz[|W;43�����Z���!����IJZUFy�N���F/�b�Z��sZ���w��B<��#O�?e�/���koO�3mH���2<dXNWv�>���/\z@ʒɧ���w�P��g���g�@�]^��Ik�\��C��
��hم��
�.��ߥ�c
z����!�ڳ�nna
��ռ����s6^���r��(A��E>����&ÉX��A�an��*�V�}���Na�ӓ]�����+���K��>���sY��I�!")O�>� (1	MJ-V�
Y}��Ͻt�j�A��{B�������P��Ե��Kq�Z�?d�f*G��ӌ��[m�n)}�|��{�Ro�C.9ŗ=���7�L��B�� �Q��M��0uۧT���}�32��My%a��x4_U:۶�VK�f;�l�E<��$�ڥ��0_�m��J�ze ,�@rr� d��+|��L������}���v$ahO�-�V��u�
k�y�Tw���lq�8F�o���6��Y�B ����w��m�1��������BӇP�4�M�OO���D�A)��Ji����I��e��Q�}��R���8�ָjޅ`�ci�
R�a�	�A�l;��&�T2��!<��{�.$q���VȤ���Ut�!��mV�M�W�SF谟8�Em�z�-�[�d_��qd+��~+	Z��F��u���$|��$�\�z��"���G2)�����&�����*�W`�t��F͎�ڮ4�>�.�����n���R�
�?���p�ף�Q���� �B�6��.Ha�Y�m�u�1���в����>�ը ��L~�ON x!J��\}��Mp���fS�q�S1G���r��� W/As� l1��Ώ����~��`�#j;ߑ޷�`{��팥9ז�����H�j!S�>t�u���	��+�Tx�7��+�9�x��U������c�&o�l;��a����OP^$���\����p}��ѱ���6���RffH~[z���F�	h�6������	���w�$�m�!Oz�Aś�� � ��4�0�-~?�� ̓iP��W��]�_��<{�Kt�*��W��%V.A�� �%n\���j��Y��V	���s�G=�t���|�'8�k�P&2���'�8��h6���A��=n���Pl}��OB�Ĩ/����M(�s�J�Be?xaQJ*��sp����~Q#�b��C.���D�ySy0���_ʗ���*v����t�~h2\�	P�S�#�-6'b7�GxB�����7+�f���R �R��8%Es��1���	N`�g�1[��\�e9�DID�;���� �)�=���w�:�m��F��}M�0ˆeo���C5��K�9�������þ�����Y�.��cܐZ������T����GpXHB�����*e�p��(���8!�O��0a�bm��Y(��
n�c�~;��]^h}�p�G��h�MR��*R����~�'HS�I#P�߀��Q5�3�E/3%��'���`���
�?#��d��,���i���tZ��y�P6kQ!f�{��/����HYUhbE��C��`�D��|�{%Br3W�-�XJ1P�<Ьr)BY��]�x<_�~������x!ec�ϸ���#��P���Abռ%aS8/��M#�J�Y������g�gd�ײ�m�_/��KI�L�����\M���M�^�ąS���4�(���;��n���
Q(7�b���4��"�x5������	��8����x����
[�����N��.�&�����B�(#.C�R�b���f2��ː����TI[�2�I|�M��\M��YVt���6ٍV%�ŗ�B{h�/ө��]�H�DD���9ړB�׻����{s�b!]H�	�H[!D�����$<+��u��3�Orc\��{��7rK��@��v��+�N��8��1����4�K� �*]`45�1,+ �D��JQ��:����M���]�nacř5�����h�������/'� #FU �wM;'�PE`��\�1E?�g�Lm����6�����|m�k���Z�2O�P���H�)u�R%c��M�lY���M&cܔl>��W�vMR�jx�����&�,>ss2��0�
84L���S����
O�o�tc��Y��op���)�
��L�f��i-��͇���HR�Ҿ�0��5��O/��T�.(!�W��VYQ�qS�Dm��MnmV,Fj�����k@����);?�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+3S��2�/]8�팘If��O��T�\K�h����i��'!�L�o��/m��$��M���MG{	����M�^n Э*��K!��,
5��#~!�Ut[�yϬ���2���m���M�¹R�b�޷�!�M����(2���9rւ����j�H��Q���	�A�n'*����#3&��b��L��G�Z���[I��qi�P�f�RK`��� ����L��9�}";�L^�Y*gQ�o��Lᇦ�X�i�Wm�Z
YN�4��y+)��פ�z,�Zg4���O-[�	B�ަ�+�~F�a�B���{ƫ���"�������ܔ�c��n\�|���w�����)�̧��GbI0�	��k���(�p-�Qt����Co, hG��p`�?c���G��$
�E���vcj`)k@Z��t�`�E�4��e��n!�Z��Jڴ�$�B)��ҽ{�W���t����?�_4��ľ�)�i�ZIi!T^M��f&��e*y��_�m������d��ː�^��ETGoq�����:u;4�P�:Nm��_
�m����7��I�79�5�-�b��aD,
|v�Ip�{�,˩��_%�1����\/\"Ҵ���g��� $����G�c)�F�H�S���6�����R�n0�l�W��\��kXq�V�ƹ�F�a;��l�����7�цO��
�X����'�R/�P�c;��K�v�7��(�we��Kl�Qe�;�[�Mh�������5��H�$�$-��Zx����5��$U���u��g~d�o��x��tb`�G#�b���nJ{��>���2��-Ru`�$��ʺ˴	3���*m@���O��܅#âέ/&.%���a�;A%�k�i��9��zr	���b��7�Ĺѓ����1��$���)B��%�5�/̸#��X��a{�+�A~��?E�%��+Ы�b�
����U���i�G��qcn�M	�k�	c�΂ui#�`��h%��S�����M�R��u;TȜ����G�L�K���ln�ʧWxuL �����z�,(��G�F˘rиua�?�I�k����/���S�}A��{X'���[�\��������t~��QOv�:�QIv�j�aO�w��x8�WY��d4��VeG�!R��m�Ab�f}>'���F�O�r�9�q�G���*l:܉�����ʄ�ڒ�rK]Әu��-��>j�z�������C!C6��`�X����gB�Q�;Y�4�m@
I��� ��������-��	Q�(áWب��/�Rp�M$�94�8����na������q���m��k
C��! �pz{��7���V���){>/FU
�����wK5_��w7�e��+�Dac��0� ����ё�b�����$��B�m��r��4�JC�s��շ����%2�}��G��@�����V7	��#3����c�Hd��خ�)]��?���jלp��X�ʦ��'��ɥ��I��f�_���9��^3o@zs��y~ �1���Ȑ+�l��`�q��䕉ǋ�@�X�i8�h��r޼{�!!�\�G��Q���2���^�;��ČnOԞ��m�������;���zء��ޕ[��ۆn`�+��"��L�ɻh{����řȥ�
�`t��zvY�Q=�?B��?��/�{}�ÉS�u�"|x�8�$Jo�.���15�d�N�K1~����M�����&��i�NI^��?��9��9�&W�����w��/'LH����s�UZ�	��t�U���~��Y�i�m��[G������}&���񛦄��;���-,��>ݰ7-�>�x������ym��
�J��!�����?`�"pyc��E�赘�ļM���<w列�`׋�-�d�B۬�>��-A�k��5W������{�">s�'6��#�i*�`�-F-�6���ϱ�.u�:a<F|=���𺵒>CkG�����������[��ǯ�������;�������T�m~�d:;�⼧�W[�f�vc��I"����oVN6#/�gV���%Y(��g/���#��En�'o�T0\�b�E����b��D�����D!��y�%�{�%�G
�"!1<�:
�|}��7�?b�&�Vs�Hm]�$�X�; ��[D|6���(�N�c׆b�ηڢ�C��d��f���u�4����p^�TL{���Y��}؆B�f�UU��DI��[j�8ϧ�G]���4�.�oH8��M_b#�N�p��W���U�N|_ʒYқ��G�`��x{�6�g�o��G���[��N�;��E �37�J o��Z6v(ڒg�n2�	u��}��H2@������ j�ʗ00E�*�7���9d;Qc]�թ�p�;�6 ��DT.�-~	eF��&U�EF�H�A�� �(ٗ���.(�Z��3�g�H����Z�҉�?��1����Q��Gf��|��7q�B$eN+_�9oQgFx��{��wK���sY٨����z0p���\�^#f�n�/!���UA��(O�^�&��]��=��=i*H��?APȟ~r\�6{\
�%��K����+��Y��3l�ɶ�/<��\q����M�7`��MhHR+�s^��N�n��g��Rw�cm��Ó�^�_���}f[6�Ǿ�3O�� �zLYU7p�Y��Ȧd钆=~��F	�%]l�1�ueH!k�W��XrdG��B���j���>+e������oL9�3|��L����[Bw���ѿ�����$ݺkG�i7o뿝T��kΩ�(ӝ;��d5���?�������x�����]�
{c�Z	��G�ʏZt(�<�Zh
 im�Us#�{&�����fq�9Ā��3{L]n�������h�$��1�¾u�x6��Q^����Cbaw�FC��](�6�G���,�p�Qd���7�9� �]��H�`|[��~%������� .��g�V.�U�a�
y���9H悫��p�&i���p�~�~�v��ty-�4�� d���}��8e��ʒ�ؒ��ʝ�U��<"�X��[T�a;��a��l,�Q�5�w �݊�i���&�<���t8��2v�
n+�T_�@*V�M]�lO�����D׃��~�$��D	�L�+��Ej\�{��9�'���i1U��8�tx�&K!A�Ux��:<"�R�	�s�*�[�I��%\���^��藚Я�?t�n�L�Ȝj�@��m�e^�X���l����ϼ�ӽ���V�v�+�[��]�-Hl[T�7W��[���w��d���k}Q�E�7s�a��.�u���Kxj`��xpLe
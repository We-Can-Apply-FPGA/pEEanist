��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�
#�i�MS��Q�
<B
�t?{�^�z����$�����Yp�Z	��O@�/iO۸�3�����p�`��#���+�B�&��Tf�O�}�li��x������2��c$����<Ԡ'��Hb&�[�q8غAC
f������8��]vʝu����@���-@�0{o>����;��9���1!(�g���?�
C9
e�Y�[� y���Ts���b��Qu
�;τMk9'i�=���h���\='��c��+����墍�n:<��UN0��k��<j�[�ȋ#+a�ݨ���Y�z�cc�PK�2�@ɭ�~�W̰l�+C�j��-o]6��|p3����8 �Hl�>���@c����h��^T���v&������C�s.kUCu����r�_ev�C��=��'y�N|�j��Mw���G�#�y�R��ӵ`�pbx:�I������� �\������a��U�{�p<�럞�uG^�/�:|�/,ϽǸo�H��7%!2��X�N$G����Gg�n,b�c���.T�2��Yn��r��e�GM���h�`d"��?yxI����*�Y�q��(5����
JZ�g�g�m!�$|���Z��CF�T�E�r�*���J�l�T��=w_pH?��K�f�@�#��<��G��Q��,���D�/���b�%��p���"�٠����<ۙ�C�����}�;�h�s�� ��;����5�N^�H.7��޼b�<ⸯ��p~1��c)˼��q���w�Ô�c���7��R��i�\����l��@l�iBB�\e�a౜��������8�������� 2w����~/�H!��'��{��1ؼ�姤���óϳI���2���.�`�����"���n<�x��|i�Z��+����S�ͬN�.1n�s���� z�tN|�%SVԕ�]G��hIU���xd��������o��ʀ�6s��
j�/%��$#���d����ې�2��$ę�WLpuė}�V�^ڇ=+!�1�
�:l����*��.Q[too��ѹ�hP��Դ�Z~4�xe;bS����sɕ���5J|8����ʣ�ZAC�2��rI�zO���mw~��$2[����?�I�s=|�c��K�.Y'�j��C��i$����"\�$T�x,���5ҼYP��E�S1����s�}d�]=Q[@$7��zM��#T�,I��R��v��c�Qs�b�Ǎ�����U��b��(n+�	����T@�f9�>�r<���NvX��p *(>��\=����m'�z���9TE#x)�!��[���:6B�����	�u�����v��=3�ox
��p=�%FD�u��0B,�Y�S���xOskR�T\�Jڣ��sA��L��N�ydg��Q%Zd5!n�׈��ES`e@k���N0��S���U��}G����h�i_����N�:�y��n�>���q
����6@ʇ'4��;��b�$o;�I�Dg8�x�X	���4�k�z'�H�q��W���*�'8��Ԓ-��+�Z���ִ���\J�󃀨0�k��e��ҿ�����4�lm|`B`�/�bQ8�y�wm�aS�E��)B+����������ﹶ��7�f-�Ԛ3���#�n%���hT��������4�b­_��wq��zff�T��c��A�6*֝΢6��/:�e6l��˧�F�R�x�ź��YGG�:��8�/���vm���וH�� ���	�}��ܱ�f�\�0Qqx&v�{�up`�e��V�������vM���G�3M�cވ��l�:�����q:�2 �cg.��<��u�n𴁁����JɃ��K���� ��eρ�P2anr
�G�Qz�wI�1mǐU�`
]<��-|��	��Ȱ �]{�Ѳ �ix���/��m��(쳨��QC�TRr�r3�O�T�9z����u:t8���-��G޵��F��%C��*|�quߘ_5)�A*�w%�(����i_��5!�ǝb<=�������#�ζҨʁ���Иȗv)m�O�+��Xb=Q� �ˣ<��ݦ��H�/}15=J������O����Bg��F{I�������#��_A�	�բ��v��>n*���s��\�����*��lRo4���X�	Y�(A���u�ا1��a���2	Zx�6�q}z��곍aɗ�j��Ķ�uq�]��q��6��0 ��7�JUf�v��)���[�	Y}�"�$���fת�X�QfΨ��Ɖ`����:BK+�	V��b��S���m'"�xQ����G��U@B~������.����jW��g�u����Ƌ�wA���>ȫ�����a�����>��]������S�_�L��%L���I$s���Ѫ�y/�C/�\�H�"w��Tp��qu3/��2�j#���*+�־+\\ ��W {�)䮍-E1�dаq&t�K��������q��Y�
Ӌں�����QnC�<��N+pn�~=�=���P�a��jD5e>y�j���
�D��mQeN�uH/mh��J��.�L��r�xVet&�I5�yI�h�����T���OTQ�3}�-wI������/r�ľ�P�o=�mv�p�ʙ�`��9Gm�Wݒ�t�i��g���	��7�P���=����m5%x^�=}�����k��'��˞��ˡ30������x��ێ�E���T!��و��#걘�w�y	���tˁ4�^��w���c����q��.���d�����=�9��%����VO��\2��U��C1QŁS��bT��EV�f�y�>"s�"	��AZ���.�̟��	��U��G�c��(6��%�s�O��rAH+�3]0�8�zF-��B̽�ݟ�{`�[�_9(���ġ�}��tG��*,�������y���?]�IR�㮓�>�i=����I���}*I��
�6��z|o��4*���v�<�M���a�����J�T;C�9�7=ڈ���b���U���*^��H_~ݳA.4�zAO�o���H]wga�=[��rm$����4Eî:�^X�\Y����l.$�廍1�"m��:y Ŕ�3�rз����돮zۑv>���O�C�j�)�g,4�E��Ҁ~�o�pQ�����R��u�����  ���g2F$�U�����.���*]ݿF\�5(�9���ޟ���錁��.�6��޷��'W,���5)�[��9!3q�[I�Q��6�^~=y�����!K�!��}���n#�w��d�EA��O(���/�V���+�+�^{�B�\	�7M�h�u�V3��M��M_%�﮹R��{[��fY����������3�Ğ{Jf��%��y�(`��A�S�i
��oI�D��;�����V;U��!����!�gq�OJ-���f3�9�G����<panAR����Y.st�{KB(��@e��k�@8@�M���a~g��Cwϥ�Ls4�X�q�{bf��a��&����Zp�^{�HWb��I�V�3ͺ�+O@�d=�	����Q����8nǮ�u�!���swԋ�Yl��'�i@�ʙ$U`*u.�Av���FZ�Z`8Y�zJ�7�����S]�J	�|��>�Ɓ-߭�Rj�p�c��8�-CjЭ8��hW����]b���q�����v,�����|D)?��7hE�g���i0� u����-�!Ԅ"4��Πo+\��D�����!���J;LUF�, ����o�$�M����5�<Jk27� Q�)펎I/P��on�&c~Nw~��/�:��Yd�o	����O��㉋4���~{��!n>|Qb�]Z���(��V.�].ep��7�Ё5�K^5�Q�=OJ��z!V�<\�Q��Ψ��%K�㨣�;��y���Hi �9�1d�op/t��`�M�(�*�m��r��ހ=��=�����?�hV��az:[�7S�%(+&�_k�"!������6�]���7��݉i������|r���j+�{��l��"�-;��� �ᘾR����ҡѶ?�b́��J;�,=Ӳk����MՕ�i2�M+`�0M�e�=�(<�%��X�gz�m&(�%�Eqh�S�F�弯�M�c��L�>��r�\�θ-dLU�R�ڳ=�u�}�'�n�2���q��@���k���lAQc��TvU��D��J��"Vwhnq8�|�m�����{��z�S~{+�!E�Di5�E-��(;�5W2���Ǥeߛ��k"�@��dsdb�f�,�V��X�����NI�z=�w�-Ph�r�%0:�UTjO��W���cHiNh|I���%�r�~2�"���,�l��	V#��#���%$�wY�4��RȤC�-��q���'�����dCcaBP�̩�~\��}l��6۳�]��d�5ur��Q��?�O���m�%�d�ZP��d���Y���M`(�b�>��|P�S��ե�8L�l�K�p�^��.{��+�66|p�N��ӭ�+~�ڙ��l�իg~�Y��(D�Ԭ���-�	$t���U%��zN#ƵѤM���bay1��ᑄ{}��X$,���/�VRF���9��Tҕ�_#~)�q+�����c��$"Qap���e%�T��f�o��O������,8Ê��O,��g
� ���L�}�k�7�QF��46@i�$����C/؞���b7��>���Dh^��
�Q�F�3��-�M���qr�l B�n��c(�������Xx���с���D=�����<1zs��H�y��Y*X�+N��#O��i�Z����!��(��M�h���8�]a\�;1�U�����	�w���}�p��F�l���|x��ݕv�0����VDCo4?`�Eqkj���\���`  ��xm�;�+��Ai0�F���P_7m0H#�ڼd$�G��n�l���o�Q�����6��9q���ɯ��Z�F{y�]J��VO#��W@�?�J���E**���:���4��!w+�X����ޞ���5Jn�.X@�"["�g��1}J�{�9������T�|�Pc��J�S����!����b�L��b��B.���Ī�C�n��m7K!����{9��w�?�y�t�W|=XݻA��$�!��es�w�"��1�}��f�mibK�xZ��)�Gy��ܑIq²�D�7�}	0gSh{d��xo��̽/�S5��!6�&�#;9�������2.��l�7�1Q���X�XQ�º���SEP�h�Wpo�\�`���M0��]Z�����X��#f\��k��C	��'�Щ��FIE�l4dAJ)���)[m�(vC䬟����`�!=�� �|�ɯ;���"y��w��V��f��9���:rR}od�KR�Ze��B)���I?e:���9*HH�:�����~'����{��@�� \J���~��я� �B��ß��	�n�!��%�qG4X�?ߠQ�k��IVH��?/���@�F��B��m�F�@T<>�6FO�Q��5n��?���y�	��՘8�%��0��4��y���=�$�Ds�v���,�0�鹮,��M)��^���tD0�}��!��K�E]��#e5����:�����oR�%���A���茶d(6�ǆW�$<|��к�w�ѾX�)b
���w�f���*�o_�͗`d_�t6Ν;��������f4L��2�NI7��Y����1E��������Kj}���1�@��F�L�[[g(I�rk:��7[t���ҼJ�ǻ%%��hA�; e�v���S�7i�'g�oA��o![$%h�UWO�O&�ze�▔�2��|W��������޻|���J40e%��E.ϖ,U�QU���ҧ���*v0�&��bt�F��8G��8���Z��󭏣����,`�	�`aC���L�5�mW7����� �����H!��ҥ�@��-�
A����&4��,�tH;8B��,`��~��"��M�;�%�V&G9����8.^�c����x�����z�Tl��Q6�p�z��#�k��߿6���F��;�K؆�\�AЀÂh�8~���TЭՊ��J�]>@��QW�_��f�����q۞��n����������� �<
�e���U� W}��2���R�@+�N2w]�Fl%�|K���ٙ��G�|��
�Do��0:`o�Svcs�ѱ�����`P1��}]���{my�_��Zx�;�C��	'1i}�����h�\����r�М�'�$���K�R���ˁu�i#�&�2�O��oCsYu���^0�GI�?�B�ޅ�J���&J���MZAW��	G}w�kvȘ���C��㭣�Q����pB˷K_�1v_C��\2_<���9�B�1�:y���	~�(+�Э8�ظ{W���qh�;��X�Ǣiu�$G���?�qˉ8R�䊧�r���䍋��=Rw��Tܩ���P%@g*�����b�K�T��ZQ|(ۑ����Jk�X�5I�wh�P��xH�]�;������0:�ú��/�/��Fuls��.1�U�"��k��G]�H �kr�D�>8�|����nE��؜��_��b��0mN��^_w��\Y�}Y(ͤ>��o~���Q!$��oH�߽7�8�P쾊�<�_r��a�����"f�$�hr��ώ�y��Q"�w�r��b�v ��u9.���b�N�|t��x�}��93��w�#�$H4�t�"Di��hs.��2�M�H$��P5��r�Է�Ϻ5`&����A7<���'��޿Z�,���X �_����uXU�L�m���� �R���F���K��>Cr�}�!HW\��_����f�q�t�o���8ΉO�{B�Ѓ�zď���,���	ln��oO�4�@Gˣ�J��J<�Ӊ2]������f�E�`l��N����)Ύ2+rX��"�#N+H�k�f��"xW����]�e����s����cэp�9��=a�P�=�_�X �K��H��I�Qi�����sz�jk���Ҏ�T������*������P��|cY=��͝�'�{�L�D~V�d��y�f.�� ������b��+��GU�~���MM���l����6�緸W!%_�|"�5�gi���<�[c#Ah�	�%�)�!�?�w�i�;�'Mn�R�(%d6��`�C�4v�r�+h�F�!V���d���3%����9�d�@�ؚ}��w{���~�p��K\[��O��l���^�&e�Y
��,�@���(�����٢=�05n���x��L�V�qi|Q����iF����¡=p ��m��؍���WE�j9Q���S��c_#��!��Of\H?�rM�w$厬A���(���tM��=m��U����G�(�o^<\�o���S~�R����¦iF	�$���g��R� AFs���~������{f�)�WRGL�r8ad�o9օ��;�2��ʰT*ņo/��N��	���GEI�����%�K�yIw�nr�)�q�P(��G�7��̌��'�L�G,V���e6�@��$�h�M���K4�r3�4;����,��,�c]ɼ٪��|x�t��d��6����=�"@��]��E�����R>���)T;��
�NG�����&S�(�I���h��6ǣ��D����hC)y�Ԃ�3���`�e6{�`?������p����?#ј�t���fB�6��c�}w��{�#�H�����Y�Ym~�VP�56� ]'�R5J�<𵚴� {?��5��Z1?5�&K� �K��%ÿw�bŎ�Aے{�;����UDx[�/2�)
��p�z�Q>z\Y�����p2�J�㫬|�Ha���~�"�F!_�`J�T��e�'t�[�|/B���09�T�H�����@���+;faS�k޶�����#2���z��-	�9U�:y���w�Ssn��R{u"���5M����U���������S�M*zn�^,+"��`��&�z�$,�dܼ��J��<^�4��J�����r���"�l�A��3U;�o2�_���Ri<�O�q11=�94`;�i��q�X���˧a��Z������N�Ӝ���(��Mn�'6r�=a]���&:v	6��V���}��kG;�$;��>�%" �0��|��B����+���2|6sql ����>96 �h$ ��C�^^�G�AS�j�lՂ�b�b�e=v��F4�zyA8�v�kxX���Ef�%����Fd��x
/0��`��6\?�~ dJ��X�)r�4�C&�h^}��<`�����RlCw�q�'gԨ���"�����7">�mΟK0CC�t��V�'���%���A��q??�O��@�E��52����%U���$�ه^��U��٠ʽ����`�؋��x@��连FM�<���X�)��uۙ^R��}������[~�4jН|g��
)�͞4Z��4hR}��M\&
1dx,��9�z��w�����F�(֑�m�������.��O�I���.��z�h�P�XA�~h��ھp�	'���]�gy�J{�����lcuKL�w���;�
T��)��cQ�<���.0�VԈ7����5�%s\&+��ִ�"���Y����{��FL�ʜ	
%4�0G�F���XYn�e$N�	�CS�x�Ӎo�2�l��om-�J�^�<�@ؐ�Lc�-��+�i^�'�:
f��뫽H9uFXk�,�[Z�?+����m�?fM���LNɐAF�H��� ���?�إ�]��$Y���:vZdң�*��x`�cL���n��<	&�z�$��`Fy��$<�GD�,���B��Ϸ������%!�h�I.��*� pg�_�M�w �?�N�m�\qh���D=�,���Q�WE��.q�4�Ja5�.�+M?;��?f��������S���Wg�k.��,]�MDf��(H�1�[�WZ�K�R��_��k�����O,����d2���D������)���I[��듹.��ސ�a�Ś�L�;w&� �Z2qVQ�b�Q4��6�m��D!�A��Oґ��@S�h�%����E�����/����o�ڡ#r� C��(o�_\>-ARC�����l�[jr�.�ao<(�>W��:�d-MM��9�L�W���;2��,'�d� �j�C��a�{��������1�]Jyizr>UO�� �z1��Z�x?��{:7�uq��9�Hh��w��9�����C�l$3���4
���߁�m��96�T�t���ܕi_}r�}�Qx����ңą���T�ۚg�{�[�I�l�����G߮A��6����x��n��*�ԕf�xfp��ɷcu�yy�ڥ�9C��q�}2G���v��
�&��PV�����Z	�L������s�g�4�K�����7���qJmf\��'�Y�Rfd�2�!/;,���Jpb�d%�:ζ��Aܐ�*��FZ���GY�J��K�K����H�^b?�4�[��/��@��k�(��k1ܦ��ϡ�F%�.��q�n��-��`�A������A��&��<�R�!1��D�=A6tO?7aOd��n�I�eji�xa������gW�(.�b�=j��N�ݻEc���c��4�n�>C�aY�^}�8Ncޭ��X��[d�!,#A}�R\މ>dl���x��h�:�W��ri�V*w�i��^���)��ƽ8w :�b�xw�W�
��!�l�ib{�U����T�@�&7��HrN�k.�4~|���1<8���q~-��*b���Χ� ��R*��v3Tes���^.r���X�
�d��B��ɑwY�J��yiЦ�ķ�	�C7��9� ��ƕY��~�p�� �k��N����鎐��D��R������^�m���[��dE�'h�2H��4����"�9��t�uYذ����mKK�(���M��ѱe��+��z�B������Q?C�G��aOmji��N�v'TR
;���:�Y�wi����'`vl�z���ںz�d�H�)*�������X�$��h�9�C�]�{�F ^d0�O��`r�-O"�O�k�m��B|�a����lt)�����t��d��HӨԓQy�J���%�̑����N0����2�6��ĘQ����Q��qYȣ���+�r�=�zV_[4�1]�X�w	U'q��]w�)�@�pE]3��?*�k��D<��}r���ZޙAR�SwF�cL�#��>�o�P5+_�AD���K=��#� ��gA�>x.��7�9��kc@g,]+���e��o2��j�r#T������ϲ�ц?���� ��j[@m�u>�i�{��<����Č�K;�~�Ƹ!�Uzυ�_�!��i�y�Bz�a�mq.�л�A� l�62���u���#.z�]ݩ`L���M���f�:�,�o�
�����y�|ָD�	Fދ�ƟP�5������Q���&
���ʯ�N� J��U6�շ�<�;��J"!�O�zu�+�u�8�t
�r���ϣu���<}6-��O5��O��Ȏ�o|0�1�1��eZ�oxp]�`��rm3.�A�5[�7�y�.�%-x+��]��*����k��ߎ|�����v�?m��a���|ܭG2T��v?��4i�V#͋���a|����!eY��#���+��>=P��NT?<����bۍ�G2�y5� �l؉L!�H�T"̇��&������r�0�a�M�x�L���V�$�>1�r
�Rk-��4���1FT���u哃x��ø��OxU�u8:Ӂ�t����F���2�aY�t���e֪��&fta��l���hY��?<�V���f{5��?�B$ܶ���1ECʃ�rb�Q��D0>��������Zg[p�7&H�%�*ʴ:t�KF�"�����&�37r�A���<��/�|�����$�;�s�s�$:���D�C�+�$������tJ�=�7>*�Y�`�r�n���j��T�r.���M1��V���;�����]5/	g�l��I��p��E�5�m�}~��QF�����(���1{3qm��J����e��O�2pHT�%@�G
]��Z���;����!E�9�����C�����M̓j�J����)�d�koi�Lٔ��q&�b�B4Y΃+#�)x�]?���ʆ��Q�ӧ>(��M��/���Ai8��h�`������e�V�#�r�L��y�ڑ��]��Z�ɸ&�L�8�|M�'��HL�Sc�B�>_��C1�?$��Fn��6,�
J���W}��Ғ{w���H�6��<I�D�m�J5$�h�5���l�l����a�22aP8 ��������O�_|��Y3��)���B�gY�82���0��$�!4
����I�t�i��� :{O`@�@I�Y���?ֳ�SG!�9�V��U���pX�~y?تG�a��סf7�p��ej�uE��I��9H�4"���l�cؠa#����$F�>"�W�a�AW��	}8�<�<�d��ϔ�;��H^l;�G����e"�hO ���2U黣@
R�#y���)�aϕ�?���JG�+�7\�.*�hfPK���L��g5��k�a��ӚOχ�L����Z��1c�(Un������_��L��a�]#�s���xNR�;�����i��PM�&;��������ߛ�284�}CI@e��x��\Q�B��1kr���Dsٴ�ظ�i�l�e��un�w^1<�to~���(�?�4u���_����W��YU$ȐN��it��<���V�. [#8��]���:�����]��e�+�C�������ע�f7O7�e�n�I�W�]�]R�<�M�L�8n��C��)�/�w����!~R�a�(�QDB?�Z$4���!�����u��<�\ u)��$�2c��#�Ҥ��������:3�.)5���<#9ƪ2v����^��a�cK���rt&�Yqzc|s&t�-7��-�M�Ip����AY��m8>�,`�6E��L�<o��<h�t�=�D��s��To��w�n�yJ�#��%�h8�1U�jYϐn�ol���7�ЅT>�;m�Ę$r_�O�#+�}ȰGO�g3F�]�d��\��aI	�h
q��C��c�C��հџUU֚$~oG���9�����dX�J޴'2/(�C�TO�{�Թ�M�N�s;��6��G�*A}IUJ��LL3�F�A)\8?�]q M�1�Ƶ�"���c/�w1����� ���
m��T�w��L|�,��7��4ƅ��Ԛ\��xL��s�`��:�^�4/1�N��n����a��)B�ek��7d���7.+�>����%c��P�'O�� �c�� �F�gg�Ǝx��L��f�=aTŶ��lH+����mNu*����-�3^�۴bT��`p��v����>Ta�j��}�;<R:�`.6��ێ9u��^V�OmF'��A4s%,�fK� �H���.�^,v��@M��mjTyA�Ȉ_�e�߾X�`-2|�~���yI�gE2���4J~�'�+���R"�W����h/(�FEXėv���!�QGM�_��Շ#���鰙����n���&�J5��,� H��}��*�i+����<E���ύk�ГHoR��*�clG0ېf�M�2u�q,~Iҽ���'�歊�س��^q��zSS�n���������{ۀ�����I�<� ��*���ܺ7���1�Pz��I�3ImW��˽�[�@e*�|�5s�[��C��8&�vgA%��!�| ��Pܐ�����*����>_qs�Ձ�dhΐZ��t�N6���aI�*�a*�է�6,�
7�XD�uA�x����m�(X�b I��g�5�v9����~�_a�G|چ���9�З����vg��[�)F-�<���O��:�RMʶ�+}WK�>O�B����W$���
?S[1����N��j�r��ɰ[�!�2�B:�	e��p\�e>����8�,�E��|�Q�k�-M<b��Q���|��M�L���+�4��nw&��ҷ���6L?h����҂Ym��&;s8�*�s/x�a;K������M��ы]p�Z��dF>G��' �~O�̵)5�!j��2b��ϴH���;.P4Eǿ	~���w���[�]A\]��������D�{��*BS/
�����䬗��j���g���P�)���5��!���{������(��<�F!w��y�����,��ΡȈ�G�E3�q�G�o7nCi�n,����<�5J
�O����i����Xn�:�4;YB&�ìEF^�C�Ln�i
n)t4R'�^��s�V9�t�xL;��zy���=2w�3ĪU��[�s����۫|D�M�(D��З�)	fE�t����FԞ�V����1�A���b�W�Q���,�_D)1�ݐ�ߣ@���?cn�q)ȥy֖�@��"�l5nM�ͤ�76��V^�4�2��,�f�G�6o܈�iUٺ�fK�Y�RX\��
ۘX�I���@�������Y'�(�0�u���V�� ����`;�_<��7�dIB���%�9hjh���&$V �z/4|��[y�<�^Ǔ�"ԝř�i�z]��*����{�6K`O�6�b
�Ye�1��t����2Sk}p��Ґ�4}Z���۳��AMA���Յ�@�7:+�֟uiK�j��K�%%�L������F�*�&��FaI"�`"2���,�[�,���	��x�|m��ӒJ̨BqȞ��O �X���G���0��U��[4>Òߞ��#�����c�M�gQ���t�N6���nnY�+,��#ӇfG�c�1���b�TF9���04�-�
2ϋr������87�u�rF;|��[�lȶ{����։�Z�� v�,	�Yv�lT�ֽH�c %��ƛP%8� ���ؓ(�?�[8Fbv�,HH��p�^�ܡ�+G	_xA���M�j��ިa��F�w��x:��7�<W�*���f�LJ��5�x�
^�� 3���_]��pa�Y��o�y��_�M��2%=jS������P�]���+_m�2E�=�W&S\�%�uK���,�r��Yɑ�A�b����9Ӄ����C��B��<zÔsm=h�fHK�V�f
�����)�OaQ��%��;rG����_ˊ'�������N���$E)��`��BӍ��&ʹ-/�@��h��E��	Q51f����֩�bQb[�J�E�Ŝ�.W���֞1�0����!.������^o�nw!gȵ�G�F���gM� �a+&��4��P��C�'%9 ���
��	x�ݒP�ab��Lm#󘲃ұU���Qq��^忤���d�#_��j��lc�qi�q��,J����Լ����ܿ��S�k��=9!�0C7�cXn:r�+���@����Z������Pfi�<鰥ZD��[܎ڛd��'*
��Z�B�`�\���mrnt�.2��5�W�5�[�g(�~�暕l��P���xd	��%�#*1/�c�(z5�M��{���0��j�&_3a���s"���n�ah�W���LܙC��� U�1ra/�m"��X����>c��{���X����p#��h(R<\��t���˳�v�P=O �5Ɩw�tQJVT>��yG�o�%��"Y?�7O����Fl����EMJIQ�E0�%�oř'�3j}��o�绱�;V�ce����ĩ�v�zP�&�3k�����ܵ�rX����H �s�(ri�Z��bE'o��Fz@Z:J��i��m��!Ȓ,����ڽ�[N	b�~W�Ѹ��3�E%3�+�����Ĩ>%&d��P�×a����FyĄk����(�WHr�UŒOs���G}Z��uUb�z��׀���Hw���@����·�kΧh��T�C2�����Q2#Og++���y�^�B$@�#�BU�8�N� ���}��~�>�ѡ�;N#�c��XLL?5�η_�e��u_���/���_� ��PN���-�����hC@�)C�'s�����[�4<�p�cy�����mR%ǹ���-�+����Hꉴ��ߐ�3v E��x9,Ǐ#5.L�,�_YE.?9�u�h2���>'3=�s̷������a����.�(	�4�ܢ3 钰��Y��Pdv���l%�(Vہ��۝[o4�r�)���ͯ(݇&���0��J���U��9�&z�W�=�J��K;h/L�oym.�O��B������`���%�{�q��s�H��K6�BU����[+h����E~:�0=�r�����5��t��=�9�LƂۮ=�ϊ�O+��,�����?�&w�Rw���l�'��<�K',�/
r�p�dQ#�b]���>������(;ک�R�O% �V���=���)֭���j/�e��&׈���l��wS	^"l��q�
�2�'EO��Ő5A7���:]�y0TBFt�Zg$t�y��0�rD�P`�;C<Zy=G_�m*a��]*��$S ��E�s�e�u�����&QqsI�U�(�<]��VȨf�~��	�鶓��9V����|��I*+�1��:1:SX!,5�4A�:kP��5/V$Av��fMb[���d%�TcM;���#|X�F}��j3��U���W���|cE>�{��Hޢ,�� �<��� L Bv�{h��#v��,�/R7�C��^�9����B�7)@y��8��STkS#q2�k�����Wl��$~��k���}K&5~ǒ�gހO��Π�(ڰ�!��G�*�I�_�k0�!����/r~j���
C������2�ɁJ��$�V]0A		}�
f�SO�ɠW/1$�Ο%�����FTKmM����W��E���	^!Q��� ���R���8��%h%�W�='�l=Ý�#����!��K���?ۚ��2vg>2��.H�T�.i��]��ϊ[}�G��,DH�(Ad=3��]�/���҄V �}{hV�FRY��5��/�A�V��k#�D�|aR��>����'p,�����4n�1���0�����[��d����K�sx�Yw�?#�ru9C`` �3�����>@�]Z�+>r�m,�LJ�I�#���Y����.&M�G���u$�T�đ&׳���B'h��|[ u�/�{
���ʣ#�:&�3/��m<_\$\K�7���E� ��ѳ�ύ�&[��Q�8�{��<r�;�D�j>('��<��X@"ϨS��b�\I��~�!�=�����qq$�6n2>�-~���8�w�M��sUF
�G����NchǨ0y]�pxw��-J[��V;6��\m�r>�L���d��}���	��PG�>���i0�/��}
�.��O��ؕ�;t�۷|���ql;��v�B&b��ߺ���%z3+x��n[�y�4	���UxK'0���ƣ��5im�� �Q1�e��p!T��P���w�y~��8��iq�5Y��ϭ�"!y���20b� 8�4㸋z�,|�I�P>�W�@�;M��z���Ӛ3��r5�� �w٨p��`�A�y0$�����������TD��
�-H� �hy�鼑���no��ĈY�;���p[��Y��M�5���=B
G�X���Ғ���F��
f���;�R���`?�V�C�yՄ����6z�)�\��up��i%|h�.�4�l�3Jsk�����:����;'�0r���QF�J%���n��<�V�j[=��vkXRh0���S*��w�*��<Fi�tؐ��n�5Mj�_����?%�lp[�|W�S�:4(�0�:�n�z9��:�0�5k�x�n��K�įB4(=��o�	��@��o��>W��VP�W�b����b�ڂ?R!�j��_ϸX^�5l['���_i%`���E�B{u�x�B��~,���:��J)��N�-��z�#6/O�Zy]:����h�E��b���߼�v9�����7#;To7j�J�u��dw;V� o�u�/Y8�Z-qщ$Ez�D?��,�8���ޝ���0�/�.�<��,������kEl���ج�`Q-F�.�D�(O�x�W�A"蝞\
��6��iU�9[���R��$�N���m�9t���[n�fv$%�f3+��k�Fts��Z/p���/k��uzՌNIj�>��|N>�K��yu�����
�͖��|m�v���t�Cn ���]�-OGP2/}��.�������JRr�ړ�i�~ic�x���Z�o�LvH�����	� [>�X�q,��wCk;ϱ��֡4��T��.�m���1�6&t������������ZT���&_�%+j�S���{���;�$U��R�_@�z`z@�s"���0rV5t�o�z��N�f�r��ғ����ұ@��b}�M} ��)��W|dW�?�u��MF����UI��کb�40�\���'.��룒�*��/7]'�u�X���%n��/OVzľ}����&��$���#-��O2[�`s��(,$����I;T-��Wޑ	��W���U�+�5�Q���tϏ�Ʊ�<1�����S&�x�UP�iմ��YȂTs�°���aӋO�N�<Y�%�6�i���4����l߸_�"1%�ͅ�y�H����R�.���]��fS���M8��d�j�:b��0ov7ɴ+&�Ek`�Au��iH��\�V��OVT.Q���<c�J��̐��	���I1������#U��tFG�����d�t
gn�"���5`��W��6�����:/#/�=@x	P�e$Ӭ���)����rm��G#� �ɷ?�ɂ܎�
�-d��.����#x~�m�Oo��G����x*�~��ă����P����.��	Ȩ��t�YF��n8�Y%9-T��q���T1�,Ko��H�� ��<{���_ �<<�:/�'��d�w��}�֢�]`�2��Sk_F.9*�r��sX��h.�l�=UϜ�s����j����\�rrXc㺠�t-�a@�Lϯ��/�����#�iô9a�x����[2:��:/��a�ƴ��S���9��t�Tb�m��â����P,���5��bhx��n;A��Z<+(���3<P-��l~�}��^��8�)�5n(����%�辆8�lD��z�ֽ9��jJR���D�K�KƑ�;֋�?ֺ�P��ё�Ro�O�spڃ5�b����^�*( �YF��;-��>��Y~!��{��G��"�Q��t]xM��������0�r/i��#|��~�!��OIRM�H���2�[�FĤ5Z�.�<H|��Ike,8��'m�0S���j��@H`r#��@�&H�$4�=#���Qq�n�s\XD�&������2	�Ə�gqv�8���𿀚�!�(<k�4�1��RQy�8�^O;���{�GfA6�k�\��WSy̙;S�~�-0m�����&ӀL��~	�ݜ�Ž\+���Z
�<��=�U[����{+=�fҤ�a�9����_����!�74��oK�����8-����1qT��H�n�lr�I��n��Q!���I�����پ��W@����>SF2�J~=D�B��#�����y��u��b/hU�[)��0M|�D�v�ԈR��AQ7|t��G:�e���>Lw#Hw�\��G� �wɢ�lP7���cd�ֱ<�B���)��}�t��pFL�"��k��S�F��z���$�s����f���$���.�(^q���Ժ���sG.��Y�s��/��Ue���G�}�*�=X%MN�Mzێ@���_:d
�-��jp�dohS���;�����p���
|��I�"�I�	���#��T���Dc=00���Z,E|k%jd@,���~m���us*	��^� ���ͽ�ܥ�#�#f�k6�2� �,��*:�ɱ��R<W[��G�e�#԰Xյ�p��]"��P\I�M 9}�+�tǕ�e�fl�Fķ�	���]
���Z~7�]k�{���1��X���?�)����q\��SF�tW
���ra�1�z��o���-�����O�m,����D�r���v�{[滵�Ԇ��E7?�khk!1��̀#>!4����첲�E.���o���T�Ǘ�ZVZX#��̇Tt_Pw�>�X��I��9��B���m�}Q��좩�/5�]�� ���Hu�ʅj���C4݊�O��]�%cק9x*����ש_�6��y�=�ۼ%X2U�L���Bf�u�3~�ٟ#Y�kò�b���~L�� �<<f����oN+��"�]�̐;>�4�e5��C�t�'���ebN�*�U6Gͨ""�p<�\�v�T&+�+\K#3C �"8a'���~h%��=a��%��ʶ��W*��A�c��k���Ǻ�%��O�]@W�s�QY��=]��0��ﴄlMs5�H�̟i[x����I��!\��j@�K����y��S-�ͱ�0�'e0�tg:�f�c����5Q��1]��nϴ*p�D��I�ǅ�٢|�ϟ}�ദ"U�@q���<���#:��Jam�{A��m棈Rs"�L�JxG��x;r�^~x���!/��\V��y��f0�W<�`W~^�����Ў��r#��l�	"�����Y��6o:Q[���Gx��E$�q�I�N�x��k����U���c�`�͢s��u�Ę��Hi�CA�;pQ�=*����S&C}�@�5v�!��4(jJ�m󟋾�9�kh���g��l/�Gƿ�=o��8�nE8�i�7���x�k��uG�Z;9�������J���!��<�gjxL����n!�tP��G�ֽ�݂`hJ�ջ��sd�*S�@��|�rT%�c,f�0hw���X�'��2���¾r��\Kλ�=��z�����P���`s���N^@k�nQ�}S��N͎�7��#��y�� ��CFz�y�m<�\AP�P=�_�'t�`=ڼt,o�w)����4$Q�$�BnU�q*��|�w�����bx�4�]5�}����t����Â��S�V�/���n�Ɖ�mݳq�$�+Qf��f�-��	��n�w;�2�I��̥���� �J��䗙����X涐�MX�H�E��k�0��g�������K>�Q�2y����c��[*A�py���j���ʃr c}L>:�­���dVX]#*�֗H��dtG��Ov���7�T��ɬw:Tz�A�Q<H7��S� �<�<��eg���C��K�]`�����%�.	)�t���	k����\�M� K��A��N4�-��K�m�B�,��"���	����Ú��x���eg���!M�=��u��
y	���[���Y�~�$�H>@�3�f<��[�9Ŝ#�y�S\d�޼���\56	T�"�?Yiң������\�AXp���k�Կ)�N����ˮ����ɨ�^h3�t���.��t�s���+�#���ʙ4_]�wq�=Q�5�J$�����f�Ʉ����+�h��%_�ز���A=��Hy��dSݶ?뿅��HN:����{���_��� ����������ٕ����#���94���	�B_g�N�"Yr��q�,F 1�4Bl;M~j��T�D���Ο����粖��'�d�e��{83�x@��Y#���}ּ:o�tr��W����s���QJ�)jP��$A�]r�*Lcm5����'��E�~Z�z.����`*�{m�"����(*
*fK�bW�P�m��i&q>h.XSM�i\)���I�Qʠspz�o@���j6]�Q�LF.0��)�bRшD�BG��_����}�a�)K��3	y�&��]�1��:�4���Q9���;�>L�z��.��	$dB�R�,���hm˨{��
�o=�B�Rh�Wݴ�N�d�T�C#[z�&R2*.��N%I�9�Ҭ��w�X�}�@�CL�ˈ��;#gnN��k�L��X�= ���&��^���C|Ѫ�Ƞ>�l���<����^{lO'�ۙ�u��c��Pw�����V�.��C��-���hf�@�c�p�*?I6|23�6�_VY����yy��!�[���T�fնCӒ�oщSr�'[�O��uƣ�^���[$����h
T�eя\;�s���;L�Oi�i�4����7�fss��J6L��t�\�BZ�~��� ���k��4\��y(����D����@?gW8L�7zNGH�۸=�Y���E�"�s��|�l-���h��G��u+�7�T���#��PV��*p����=�@�)Gq�����S��o\H��
f��4�M�+Q�E\��.Tc�jq*P����F�q��މ�d!9A�"H.��|�A����h�d-�^gd�'a�O��7L��	}�������t9�j������6��K�My�G�3m�;�|��9�|�H�Im���q�V��a��h�`��jUTx�4A{��M������������Їڐ�bv�]��͘L�P�H�i���w�n�ڰ'��@����d�0�tY31Pz�Qd���LN���� 3@fHFGկ��@���b��T�Ҙd��(���|@�]�٪�)e�f��*��=н5=�R��L��-v����.��s��O�J4�Q�����������Y���p_�͸�F=ͣ�޾�,��N51�,���вj����$��$MF�_m7��]&��x�7��F�åI�t���}a�b:{#�2�Y�ظ���x!������ص.f|����F�L9Zs���b�굀B
�S�f��,ܱ����h[ʥ�~J�몥��<z`�UX�/&=�/�ix�k75C���*���w�Ǧ$^Kb�c>�K�n������{�m<l���\�~G@�Q��S��G�79qQ;|�b�*����p�]Y۝��	<h��KՑ�����Y��ٷ�7�3Y���o�y�$���0�d�'�e�-_��ߝ1�/��Vs9_���!������]�d̙2o���s�U��� �2�YB�d��>p�"z0;�i���U*~���u��	�l	����B&�/��r�*>YT��,:����a�g��ô�7	W��d���ď	��Mh����89��J?
EQUazVZ��1�h�h?ɟ5>�\R(�'�J���]�dl�M@8'�b�?��7�% �>��JNv�VSWQ�j
bߙ��������ɘ:_瞅	�<��:�۶�^�fsZ��!� r����/g&���bix� �f@�-��:t:^����i#Y�{x"5:��\����p��������yJDr*�&^+���F�Z��5������b��%���E����e��������j�J=ZQ׉XH˃u-����9>y;�8U�j`��W���!^b���}C�X�7r+$���b�/s�}� V�ϝ���uQ��z��L�wg��*)�� 	�]����T�f͕N\������_$��`<��^�J�c������{�(E�]��<Ķ�3M����R~�LA����M6+k���=N��m��|QQ��]?��c���dq��;�����d�K-cp��q�]���S�@T��t��p�r%���?VT]~ԃ.�v�I:qr�}C@)5V]er��q��x�#��%�]}| ����́�L��'��9�G՘�p7I�L_8����jP������'�l����c&�����A�C䷱[aG����'B�D�x�
���2 Ky>Tύݨ*�؞����(��p_vd��}�K����y�,e�Fv��f9dC�\1����Y���E���P�i��b^/��}������@�`�A �B����y1����[�4���q5=k���=�a^�j+���%S�J�3��Hq�4ԸAW�[�����/�3�ͅf�L�'��4��%�;��/���&���|g^X�`��C�*V��*Xx0C��Z�z�c�ߟ6�R����)@�����Ku��n�qJ[���T��&/e�\`}�R�[S�ڹc�N�c���z-Fɭ`D�lH���bj�^��>���dg[���)͜���b��y�J� ���Ky�=/x��k���H}}�ń�{\3s\���3-enu���<�L���3n�*R
�R�>��X	iyʲX��9N�C+ʳ[�S�v�t�ږ� �������Nt�p�osJ��&��Ⱥ�q�g�����:��.�P�'z9�ͨH�t�r=R�2���D�+ XZ���>�3|o�^��|�H0�ou~��{1-b�uo�#R��k,�Gn��+"��F���kP��������<�faB��J� �[��2����o�3���]$>��cy����?��R��F���ҕ{��� U��~ך���Z���,���"�2���񜍔���j��J(���Q�D�h�<ãDʑQÆ^[O0�1�kI#�\�&uA2�EÒ1��j����4:k���H+8�WŸ�l�X�w}�.�:5�����>�d����A��i�9�>d��B|��k�Po��m�}�
���&���Ccw�i83��%�h��̌Jm�i?k�L�~݈��c�F{�X�x�����sݶ���`��eE��ԧ'�B h��L���LR�k�|�NV�� G\�9k�6e�m*d�9Y� ��4��(���Qd8�F�3R��o�u�hLR����B;�����$�#�RrT�Xة2L�����jS�ay�3���q�K�	����n�˝�o�1۫x�Zh=�r�L㓶�pK�֒X�d�-=ѳGA���|~#����-���2��G}���k���*'O���V�'0���Y�FIu�?�tG.�"�'�sz��l(���§s� ��+�몠]�ՋG˹�����M�P�(ˆ��yá�駄ni���d�!��ε�t����S�O�;uCp�r$�m�]T�5�~I<��	���w�J���O��(�ˎ��vs[���G��J�/�g�ƹyk�`�9�y�O-��"}$�H,k<!cֽ�ѽ��U��ÏW$�<���$>Ʊ��T 1�&�Qoȟ����V���V�3�hlE����M�L���9�<���ȃ�x�a_>����6}�V�՘��$�	qjw¾�	yW;�L�D�u���}*�>r�+��K����������0bt5w�}E]]蘫�F�x��!k��nZ�5G��^ׯ�$9j$h�T_A̺N|������sϛ�If$��jz�~d|��8	2C�*E������5E���`J(h�gx�wҚ9��wĤq���2����IGo�ܠ�U"�a��H.�:���HU�����FV��ꈷ�::���퇡|Wb��&+"�}x���cs��4C�
bl[��I�_�G��43��bo�nkSꙺP2FR"e�gm&#�uOT����:���j��P�.��i�D�ܴ=���� V�R5����Å�l&��#�mKV!-;�_�R.@�����W��yïx(�5 m�'3ƒ� �6�)�]�N6�(�L��m�^�	���q�C�����S�=>`mUK��U=cee�Z���I�8���jZ�A��E:t9bj�`7u]��=�q�;'C���q$�[܀V���N~��O��!N����g�P����~����"�8�ʯ��S��7��y���K��g���F��D�1�Me�ũ��s�m�&��*��H����S!���u�k�n�<�e.�h,�ĕ�-{�f�*`�w/�)����pp<�-Ր>�Z��A&e,,�(:㤬�`)R�q=��*pRԹjn��|��Xk!�Kb���]�#S#ڿ���h�|�
P���TF�U������aHUۏeF�c6�x�2� �Z���w������Vʤ��п�(��-f*�=�پ���4ˏ�!���Ȕz�h7�F'�V@CUy�p�f�T.�fTHk����y��T$�Ɇ�Ù$i��/��UP�&ȴ�R�	����3cW}�Q�s٣�n�ө�V���p.�1~�vP�c���Rq�Px��:��X�}=�V���k��'�z5�����2����SӼf$�,�O5�B;�:Dǧ���q�U��g������$=2��J1�k{3��4�B�B�>�;MY;�
�c,fꮪ=~����]x�}.��<�����鋻&&�킈Ġ�`�q�vdL�'ox��$l;���ί�3#Uoz��n� xEd`/�3G��l7a28X����Hj���*�,<|܆���}A;�\� �iqP?E,�f�i6�ʡ�}調�X��+֢��r"(1���Oʴ"��ҥ�DPd$.z{��7�i�#T>��A���1�:�K:���,�!��Ό��k�C�L�/���-�����3�_��Z�
�L�Jz�z-8����R�lA��
@1��
�&Y1M[��R !M��k�ʲɧ��G,��L�ʻ�Ƀ�S8G>�b�W@4)T�
n�v�g��,}�t NAJ��,F�Mrqe�,����06������(�+,Ls joG�5�"�oD�x�Re�z��027��>�7�T�5�qy'�L�V��	����p&��'U�v�����]��h��B,�>M���Q��N-x#$���[�����\mg
A�J�0jL�w$��0�[��rAv��p.vۓ��?2t"������;6��`:�v5�W��p��G���[��C����WS���uy���)�� �juٍx��9�;�E| ������sG����)��tH	:�V�=�4c'�v�Q����H���ϭq)�|��kX>��
&�N�����[,5氻���1bg�m[�1�|ו�c/#�x"}��-�ٿe�`UE�5���\��@R��Q�ZS�l'rzU�T�Xp�x����~���hCݰ-��)\�#�;ó�|z�����O �ż�����X�.��wO�^P����ę�(]��)��ڊ[��n����tVd��q��s����l�JQ,����O�rITH��U9�}z���{��ov�x�8^Huxa��j7��u/y����B���.�΁�Ԧ�
&%�&�I!�)-�$v����-+��:H��N�P�o�›`�Ȋ�����Yj�(�����A#ԆBvE��	F�3Cm�^�� ��r|���t�p#�׆���GަN1��k���n�
��f�=n}���؋l��,�Z��D�b�=+3��r]�v����d�9Oǚ� �$9aB��^�'��.&	1Ď^��M
�Q��i+<�sp��3���y�b�稌��L\��`��V�9ˣ����q_F��dѫ�)�� �x9���nI������d%�X4jyg$~���`ڂ�=F��:ֱ�S�) LbB��֛�y�<��P�u���&*o���rj^��{����0�e��$�CW�!�Z�A�������)x6�V�K�o�eXp*Jk$��x����m����g�"���pW>�Ɛ/b��﬛ڻ�p�!u��B����h ���5���gE��=aoD ���F��!`Vn��=4�N���6FtF�=H�� M���{������o�M?�qֻ��I0��}!����e�{��7�I�׈�����������xk���n��0	�I"Z,��H�i��ɖ����q6N�x�Mv
P-%������� ���U��<J�n��G��U.}��G�+��|�#SQD@�\�UP�ޢK;�T��u3y��J�֣�O��D  �$��P�_������|B�rjTδ[y�^��,���~�/�y	'���=��KjC�h��vTŻ:��Ūj��7�����4�[�ȼS��״f��{~���;U۸��,�r2�a�?0�}�m�o�Y��b�)�x5���^A���Ⱦ��H�
����DQ�wa2M8����y[��'T ��[��1i���<���07��	�}��!������3�a�Ch���+�����[Fis1鸠�9F/��W(����_���rE���[�{�h�-9詼���J��e� �?�6 �N����}8���4tfmRg���#����X�j��`�
�Bd�z|^n�_߉l*��V�?K�.�:�ݲ0Τ�<���yeAH�Y���׫d�oJ��R�wV� QlT�h��NiQ��O*Q�[_mc�?�5  ���#N1���9<���z�Ω�s��W�^b�j��F�A�o��
^�2/�A����-�ꊗB�@�{�$�f0j���ŗܥ��D{y��f�EpXXwZDYZ�։*�㩙��We�ns3�Yس$�K?�)t�/v7���g�Wn����p �����g�P��FG(Р4�K��}�d�|P�;a�;ݯ.0���d�F�暺�P���D��7A�e�1�2F��c�`��)4�P�耴f�q��R�S�'wME�1l����qx��2��	O�eʏD��R�	(>�J��<���|m��� ����/��/����U:+��УR��~1N5�K���]�4�Ɋ��%��*�@�4�l#�ڡCy��u�ϗ�p��"���$��QJ�Mp��}� M���=Tp��� ߺ�xѩ}c*@I؛���C�qϠ+-^�k�`��2�AO�-�_����/��kc~�"�Ϙ/9i =�N���qSDz���6SH���/��.�@T�&le������˜�%�SH'º��������8-��|���� ���'	���p���H�)�%�.W��C�&�ٔ;���Q6_�� �/b�?W�?�sDW�(��,	��p4�`!�(��@�:���2����a�PJ�)�]tXH�	���w�XV���h	�^[����o�LyU�++ z�rϥ������T�\�
\UŢ�9�n狈&x�xLѓ
��\�u�v2��58w/�	Æ�S'����\gC�#�T�,�'ݖ�2�rǊ�h�>��j��~5�7z�Y�?Y.P�@>."�1U��G��Z��ꝅ�'I�HD]$q�xF��Ww
8�]s`�F���_��g�	��Z��=�C��?�gW�Aqo<�f�᭸3\VJ]]a�����,���.CSQ�C�~�)�,���i��~.��np覒&��]�<zFd^�"�"��4m��A���L �������:�#7@�U\L�e����kj�?wޏ�%D)w����>p�����uI�T��X�j�F�>x�	V��}5��}Q����5�M�+�5j�=����9J�@� SC���[�/N���%��m%jJ;j����O�J�D�p���NA���:���JUf�M;�r�n�`zS,�g��xA�@����Ѱ�9I2=yy�Hs���h,1���w%���?��d;H`a��n;'���1�(�~DsM$D�%i��S���'�m�Y����C�}N��n��,�_^���3,����;1$�h��Ri�	.�r�Q�pl#e�P'��#���E��(X>s�jƔm�цi'��S�.e�Ge֩��gg���g�b��7�.��Sۦ��薪�� ŗ�jD�%run&������%���[����c3��U3�<M��63�����oty�w�ڌL�C��wk��r8��+�N�:8+��<�^���Y�������=S�˷��|��N��Y6:�ؑmwѱ�&}'	ĝ�Z�4����Q��׿�s<���2�7;���y5�1f�Mm���k0=Oر\�%S|i��?j/[ZV�k�/J"����FЉ7��~e�I���$��]��g5J��DLq��}Kџ#g�(U�����.
S[�j"�I����`� �Y;"��X�7��'H�J��?z*�r�F0�M��"��z���
C��2';� �ٰI��}n����� z__8M:V����k�a�ȳ��������Q:�?[�f��i�bt���'���>�
3��%\I��o}B��N�C�W���O7"Pi��$p5Wpf�-ku�]��w΄�J1��\Q�����uf�T�=��dW�*k� fdG���I�)�K�@�˓p?�*l�Sse	����@3�e�|Nc(�}�)}�r>*��g��`}�w	V�_���Ka�bT��֫��K͚k���|wլ�����.eMPZ�M��s�C�1�Z�
<��.E����Z�O�+�O'�4jW�I���d[&����L�G����Ͳ%��쵹�d������	�_��
L�һJ%���	���Օ��#�`�:e�.�����S����j?Ό�:�IB
 Z�,V�?�!,~U��߳����6�}��D�M�eѸT&�H��lf]��;�ل p��|S�K'��__�t�1�� �����ߴ��US!��P�L7��Z�F6HW:��	!�i�)�%���~*(����f�/1����������8�-��9�0����-R����~�O�y7���.u�7ק�S�ѩ�n~��ʲ�Jb�0p�g7D���s�|����v�0�	�I�}T>��*��C�C<!Y=�P��Mz�a�uB\Y��h�[�4�A��t��������?M��`��7*�C�,	��\iT�'����jq%�46s4����{Z��!/a;8�i:�p�F�9Y�X�&
�6}�"~���#����Gs�$��b�	�>�����gd\l=��R����c�����6A��E3���Z� �̖�cB/���@2����]C]�mHM�������͢e��AB�v��_�G߬/8G� ��g��ΰ�S�f0��g��g3
�X)[�l�)|�Ơa�<_uUĮ5a5��=>O��X�LIk�'M�.��T~|�f�$�GPq��me��!;�<��f8HJ?6,C4�ҹ;���>�s7�����T;IKNodNi�Iad�̪?��q��23��?Eq�µ��1��:/�z�sMAIq��uz �#�I�Jɸ�r�(�#.#�`}�~&��\ %��ѿ�����BB�(���Կ))����l�I��a8ma����<p馤t̪.��lR��R����'ń��q<����@qW{h)o�
��w�q�7�!:��,�B;���6O��t���s�N�{����.BsD���շ5e,�Ʒ�_&ef���%,,i��u5�{$]�L�$wmLɚ*�0��G!��e�F�x���@�}܀�)6�)��1�.�+0������b���{0m��[c�$���������nM�܈~�b�AR�`BK�rM�`��*Y"�:��1�Q�1��e|� ���&���4U�@F`���??O�4M�#�B�i��,~Hw2��7�k�σ�y70�*U��Ɔ�����%tBg�q�k��c��F��.EG2P='������'�|�Ad�Ոc��Z��=�ts�I��w��k�Ci�r�JQW$��E"������uV�p���=S# ��6��ͲU�ㆋu��ʿ�ޯ��t��5�t��ӥ	p�)gi�g=�nK��B�����#��@�A9��f<�*Ԙ;\����6�ʮG�U�FK���7�G�Yx�>/�@�֩��x@�IF�}��v��186��{F��$�B��wL-m���ɏ���A���ԑ��%�Ґ`���6sM���,%�Z��q���������4��T���-�t��1�z�Z�Aw��0��Io��T�~^n���kz�S�!?"���X��\�8���Zn\�WR�����U���	��D�
?7Ѹ��yhR�%�2T��J4/,S�M��eT
��e=�k�Ė���?7B>���V�M�I{7�e��O�`<��ɹ�P�"*�����U�>��	nUg���^��!�P�oP2��c2ЩR��Ka�k/��vD2d`���ۖۅ��{SЦ62+Ҥ��9ӇF���/���b���	R��^��C�z��!����nRah�m��J�M��}�ǻ�ܤ$�ȁYy1N�ಿ@H����_4z�ȫ�����;%$`���} ��F��V�O�g��Sr{������9���=�d�����4�Wv4�	�ġ�9դ����|���豲O���u�V.�H����j��㩖��n�F�����A$Ȓ�\��d�hgdt�@����oQ����e_N��HD$Sw;ْ�C)�m���d|�2)*�09�N�s}H%����Z��C��AŇLxei�b��C`����'R�;���\@�]�����(Yz�o��fi�ϒ�1�~�����[Ч2q�K42����j�+{s^h�^��� ��^� �8��͋�u�=F{?��W��@�63=˒�����{���4� B���o�����gF�A�IEaz�����}y��˛I����C���i`��ݡF6�xy?���U뮫GɥҨ�_E��w��7�n��0�ʗy��a_���j�4���-͐e�ԣ��t��a"�lN�Ҁ����·UpǬQ��wŃL@7{݋u��E8�o4�	՚ڶy�*�������<�g���E=��*
����S ��N��y�|�ѐn��oy<�/�9ǌ(���@d���j �
Ίp���w�r�.@V�4�c���
�_:Zbu`Wě�Fƥ�6��B�V��oq!r?�%�F��͛<����*��.>�B�ُ�T/U��^M}x����r���$	0�3�����jlo ~�m������q�\
��zr�4x��h�vR�F�����
t�^b�Qdh:%ӷ���M� � n�������`�5>�FNl��ܹ�j��1�hJ�?]oc���;j%��G�i�ko*gֹ䊰G*�9�<���$Ѡ���Q�P'8��SQ�O�/��b3Iv�R!kBp����9˼i��w\�,A���E�D&���R��S�id:�7^�C����UK��&�z�NSK�?�]��}dʌ�D�Z�J�N�+<�k$��h�hM�Y�XB���瞂��|
h�f )=v�O�5�YG���r���]i*#q�VN�6�����#�	���Qr[��!�W"���sa��	����9����ʫ�g&��4��k�4��.���l��aT���5�I�e�q<\�>ԥ�xge_'P<pf"�mj�yfr���v�0,��>� ��>���etg�-�|Y��Xנ@
�.H1V�rǵ�sSjf���T!H������f�ۋIפw=�pH$��K.���ٕ�����r��ƨA�󀀇�2���2'H�;�/j����ܻ1��f���f	�Kl��Kk�u�`�sFV/��}9�Z�o��,K���`����\���W�[�s��q�|��TJr?-2�n 9�@�ņ�9l�3��N�ȿ�M��{���J�ր�����goLl|�ʏY(��#�n��jc$���r������������ߍS��qK��<,������ ���!��9b*���� 76<���w^�j�8��F�K�L}E㝠l�����[���A���^M�6�-/�,PY�,�iΒ�|	��Ȭ�6�}yEkc��N���KV5AV�1���c�W�Y�~���~�3�.�kxg������V��I��.��(��J�pI ���[6�h7��Sc�$>$��{N9E�C�AX&����*zYcޝa�3j��i�V?X3�|X���p@u��af�iqd�����{�O�`�[��UW��J�>�4�$�B,Z�����	ckD����7��nDfs�--��G1�_M��p��|\�;z`;Yq>%� 2�tvBụ�e���r�`k��1Tڎ����L�?x�O<�|5ć�����X j0�Q�|�:���*^h\��e/�(8`h��f&g�h�^�g���0�#��,��5Kkعe�~|�1+S6�2q4�~	���ă��3�Ѯ�g�+c���>|l�0XHˋ���DɦF��'�`���)���Y�b�h5 .��#1C�s����' -���Iyz�<O+�DF�nܩx�[��"�qJ��>4�����y�W��o4�ڮgUj�r&�$!���PpC/���"5�F�u��<�8�N>H7.t�#4��x�J����� {�v���z�p]�R$%����!�����`���<"��{8�d�r���G�{-se�H�l�?3���5��9�E�������6��yV]_��n���&
XZz)��2���_łAL�n(O���|`� (��M�kk�⨨j���Hu��Q��$;�ȵ��o3~���Q���9�&;p_��R }�#����;����bZ����ADC+�F��N������Vv��})ͳ�V:�n���`��<���Tq4�Á�Ͱ�\h�S{���K���6G	�"�4m
5�n�W��h��S���G�p*��L���j�$�T�$���b�����bQ�|���D­g,'��O},��.��	v٫|J�^֩�? i
Dd���� ��F�o��e%�Q��=@�:Ok�B��c��%�ԓ8�<m��Tź������33��~� �R*-���{{��q�iA'	�Eߑ��f������dl�	@�ஸ���Ϸ��X���p,�]h�W�Վ�bD0xܷ"E�������<���Εz_l����0��<9�X���i�\ p͕`�,�{ю(���w��ikBvJ��]DPZe��]˷�Nj��իU�tĢ�p�i<�t[�VK#���g141KV	��a���YZt_Y,\�'���]s.�܀���[� �܌��e�S�#��E�R��Ah���8�E�����\������4�� ޝ�0Ғ��⬃ʰ�ĳ���صj�\~5k��,�U� ���^☓�3�^��1ĦQ��n�~.f 5o�����-�^ʜ�`xM�]b�w�\����Ļ�U���ĥ����7��(S�M�B9����ţ3x|�}J��1�՚\z��jM��C�Y ����D���HDTX��)�WD��a<��y��`D�;����qw&Jψ/zo�DD��Z5λ� ؕ��.�]�y�z�>�'�Ch"&_�^/���8 ��*����h��M~�p��ǲ!Y^���xj��mǴy+��^�X<L��dH���=[n�f<�睜<(�w��Q�����p�����ea��5��Q��H#/�M���>3��(�߉�J<hܹ���걾Znn��=�2V��ڦ�p.�͚)�9�<x�Y���V!�tb\��y'���q�_	�N��q �?ED�'�T���[K^F�0k�z��(=��}'����ɀy�_ϻ�x.��q�����ϊ6�I�`n��8�֩��l4fͶ�o�\B1T*b��ށ���f�J}|#���%�Ͱ3��dK܌r<�/����I�J�3�jꭹ�0E��t_���|OVUƉ�8�cU[�,���Q^�E�|t_��t3$M����Lr�9t�X�$[�f�8��g�
�P�I�٥n�{_aa�a���Dd�w��zw��Ghe�u��b��9�*���Ӣ�Ɨo��[��$���GVZ�?��]`��3ʪ�fo�P�ɻ7��E+?j�1!�~>!����G�P]� �b����g")Zka}i��X��4u��T��fZ���f�&�'��6��S@��]�MÖd�	:XU�� ���&�qF|����@�Bݥ��uc��$�M5RcӲ|�>��wk`riSq������&������y*�)c�����H�R~���%��WR�HV^=t���x�J2p\��σ��м��.�ҿ����S�*�Q�7����'@ G]��ٍ��:�$�la."�7?S_s��{R��|�9�iy71D"��t��b:b�jr|f�2yݱ嘛���9�����@ۡ{�? 	.�U�Z{a|2�����tOZAz�={H"��a�-�2�j�����\���p�%ll+���A��D>|7-4T5�<?�X�2���9�p�#𗞌�&^�Ɇ���Ay[8wp��V+}�`$���s�s�S�an�D�_�خ�h r��V��F�A�}�m�,���B�vU��Cys\����_�̰��U������{1u��g��H�X���x��a{>O�2o]:%�|��5�R��$����xp`GA��y#<V����8k!��̱���H��<��_5��մ#_F>�B��[�/C����eU�Ϊ�["�L�J9��6^�,F�g��K��b�ʜ�ϙ9!�@�}	���
Ō ��%J5��;�/��C��4իA�F��/�Q�SН��b2���K�ݔ�I6m��ǰ]lƫ�q���Xt��(����%�/JL��0y~�kx��J�������Z����]�*��)f�ؙ�v����bm���sϒ�"��+�3}j��Z׋���G�rF�jqB��E��u�B�СX������l! }�h��1����mB'_�G
>�^������m���P�c$%	�vJ��L�m��fvJ��S����[֢݁/J�O>��+�gn;�f�O�q?�H��!q��3l��_-�*=fr�Bir4�]���QA/+����w��F��'{�k�r%�U����~\���-��p�bBj�]!L���v��f����W�û�XU�3��.��FӅ�	.��tp��X�h���M�A[�
^�> yڝ��� ��qt��j0
��fZ݊LI���Y�c��R���
~�0������k����B�p��h�>"za���'���,^)�z�\��/���;bzp�mf��T~���8��*�g)��w��6�u�bT�%RWXR�5ӌm���(�@!�����3� ��IqLJР��Y��������(�/kp�L��ǒ��-,��nQ��7�ߛ�r|��~��	��1Op�-�.���`�B��&㼥^"���-7}���^�@ޘ��J�n��L�+Ża袚j�FOr#�����lrUȏ�Q~��H���|W�[I�����1�R�:��16E��í�����9L��1��g�7h�����'�����YRn��ܻ�+�G�?�I#�uE��ץ;ʕ�{�b?��j�z�l�tuf.�)���A��c�����s�{�s����U����\y�𰏰��6���RZ��s�2\�5i�^e�Z	AT;�q��^�>���>���(<V{�����,���W���x �)��=����G����sٻ ��Vt	C�ٯ�uJos+1����N3n���p��#غ�ލB�OQ��X����e�=ˏ��au'��y��\�HK ]]����㳑�d����ƹкX�գ��� �K!0��K}����w{? �� �u��Ai���<��g�(}��iX'���3�^�_�+ZM�HO)\���
R��1xs�C؃BL�p��8�~(��x}4�hT���&���ƌ�a�������
�a�� �o�j�f}k�/W��F�J�_��'�]�Y� �%Lt��TY���/V���̫��"��=�����UȝyO��S�t�IB�u��'��禁PO�����h�dXQ@��H<�p|!y>��ӛ_��\{����Ú�"}?�(j�Y�o�Aj�t�qq����iSr��UML�P�7^���WD�"�P����ż���U��F4 �<�+6u�{M����o��%�jńa��7S�v<'�=�~
�����k� ڕ�TR��\�~�Z��Df�����"z�x�a�����s���t�#�j��K,*��;=����RW�e��U�_>Fc��W�J	�v�yUN����,QP�d�\{:�=�I��!�y$]��� ��*��2^�QU�٣�	{IdA�\\ȟ��Կ�#�v�@.�F+%R_�������Zg��Ѵ�<��E��8�r���:Μf����\�35����x�v� ]bxʫ�N�S��֖5��ӣ2��H�(Wن+I�*�+�P�b��x��d[MT�������u���	ѷ�x;�G0&��O�|����m	�{4Ѡ�1@�!(ӹi�-`�� �����F��paAs*D ��m"��:��T�2�����1Тp����(�w���z`��I�6H_�.\	�5/�W���1:�B��{wR��U��E#%v{�\B�h��hx�g��J}����_9o���d|���̠.߁.Q/ꊋ����Ey������ �#��!��YkSԶK�7�������.�.����)���^����@7�
6�naW�����Qx�Z�toj�G.s�'\>�UN��k�I͋<k�Q�8�"Z� U��k"�e�ij h�Ds�;�V	K��޳<�o�}��F����d���zX�#p~/��qn��9�����g�oKe8y�)Nwp�y��E��ad9����ͳ�����ҘlfK��Nݚ���W�H����ê�[��|��r��=r0�ж�%�ǳ�$l�U
$N��d��́@�4�:��p� � �p�=���(��U[����n�iS���
2'�:~��
����ȡ�2R��B��|yQy���C�ѿ
sM�fq�h���s��4�!��-a�3��0P]���+�1�����^2�fO�����>��q��N���V ���y�Us9�j�%�Fp�K+?o+�=�n��c��Q���}����o��c�a�BP1�{��wAʄ�a��\�)��Ƕpys�ɯ�Sd���dmO�Y��B��m�3�|dHv�*����M��y2���)P�.�A#�1\�v�"r�����W)=Ub��	ɯ�4���H�Js��������!�E1�����[������F�)�L�@oǵ�uҾX7�AvD˘`��� �,x�8i�n�/�8�O�T���bnV1VXtqa%J�7�tUM+r��ģ��l
�	����{���| ڋN�+U����Ǧ~���8��o����ٯ�$�(+�Q(�~䅂�n/��_k9�[Ê��!�$�a��*���ׁn]��N���6�:2�V�5s�� ��%�m���R���R(���ۏ����}K��'H�t���6�R�;}q�����m��Қ�D��/PP�%���SN��N�#k�q�	m��m����o�n���|��θ����:�ⴖ�<�γ�����Z�an⦃�L��� #B�ʉ�V�O�,��Рg�!��6�f5F��UP��	m���㻀m˭%Q$�50J{��� ��|Z��:����.���.K���_a'n�E@Fd��k5J&�f[@��r35lg�()�&7>���z�a����;�s����lݭ��yLȜ���K�t(S	O��:�Ef�����`�!ֻ�1z�{9�����^G߃��CϑՍN��h�ysu�Ͳ������B�8-�����_�TqU�^��5������i/�K�������C@~(���O���5�8�~L�+�1��4�w�9l�$��7Cip�[�+qW�M��u��� �,8�
�v��n[�m������h�|D��dZ/�����=tAn�JgT�c�	�<~6�'����U��ȇֈi�F���	���1��K�ti�Q,�c�m��,�/,�@[ߣ�,�#Hb�B����F��%_��}%Q!5�������)��-1�M�p����?�� ��Y��	���4;I���sOu���<�$Hl�휗Xv�3G^�(T��e��yn|�W�x0$�
d`��� �"�.�Э��Z��qWjxp��^`�#��mw�fI�;o$�<��l����q��4@҉�H�Ё���/Y�^��e+�ɫ��6Cv&�}�.����-��i G�烙���.˂n�%�s�5�^ӌ:{k���>&�����
W�Cd�ug�O�BF@�)zW�46�lѬ���^��If�{&�����٬�&o3V�%����;m�T�D�Z�����뿮��!R��},o��L�W�w�bؕ~�.!
���l����$C�F��z���U;��aK\FS�/}op΁
�U�a��c��GW� ��6'�)	��}b��M�q�&��L|�y��ce]�qe����g���v�L^��#M�$A�D`U�r7�/�1���VZ�O
�C<��j�](2��q�Cdc)�Aހ���D�Q�X��ݏ��Hr��
�����I��~�K�@��<��O�V��)j�A�P��G��w
	"�E>����`Zs���w��=��>�
�]$]b �_��,`�B�ΜM���� ��b��У�(��iƁ�F����C����-u�� ��/�(���R�[��C&&���&%"�wK(�=�#X���\H������s	P-����6G7R���F�
�
�O)'X�֐����x�p�7�/�t]���_Ơ'�[��<X�n(��ʨ��X�7�١�qh�{�H��K�]�!Ob=Õ���Ӧ��`F-V�m�8��I��_�I9�z�;X��Z4٫݈��.N˫BL%�$�$ot�uh����oo��7O 1����:��l!-)��Z�D��������O��Xhi�_|Ǡ]�#y>br��*�a��d�舣SiՂ��}�����'����WLݘ�p���,+ﻄ��ɼZB-��p�ԕ�CI��יx���j�T�M���I�N���Gǵ���Ȅ�&T��&�7�Յ*}��wa�D�4�m��)[X��&'�������T���4T���b���B��|����&#\8w�A1�Ѣ=L�BQQ�� ��|��f����s'٤�A�*�X)��^l㻯�?��6=x�����	'�c�r��)��e�Bo�t��J;���(y�N�|�uT��w��w�x�aFP�Cȼ%���X��e����ZO�\�*���!0pK���%�9���+
2Le��@�/����Z�H���CI�x�Q��B8���σ���Mz���Z�~�D�e�aƁO�h=���3�X���rBD�~'\|a��v�.�����?Մ�c���8���g��fa�$����F����	h%���r��e��7&�g�KhS��.�)�e �h'^'[��B�����ܒ��w�jL�����Ř�K���%�����3�oCɁ���}Uy�����wcP�`uGL�w��H�Ya����r�*�Yr�3ˊ�,��t�J��A��6�B��h���e��[��4t��z�2����7��7���p6��d���m�áid���j�݅s��Q	�U�,}��V�ұ��WS������﩯��&�i �O��z�e���^���P1j�@�V���K�_r3H�҈G��o��J��	��7t򯡻b�L)�\v.���-B/�3>��hYvv��i�ƙzt�<��M��V�8��bg"E��!B���/�����0Zf~E�����ϻ�C��w}|4�ذ�ҐpA��h��o���x�v��IE�^Q������|U���Dk�к�l~	Д����q?#c����f�c
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�ؚU�Uj��_� �~2
r��nA`|~�	���11G�)&�3�;3��zb�o�$�[���!�����3�P������LXk�$�=�uze,m��I`��
�`2�:|7��H7*���haH�x���6��z4��Ċ��PgO����჉u$,=ğ�m��:`�� m�X$ɭ�}�=%�TQc@���r����.�K���(�@��
wܶ'2�6/,Jւ��Ѥ���xKYN��S��H���e�������E�������Cњ�>�6��a��H&�fXW�v��<�3�:�oc:Ŵ}�L��������E[�͔�D�����p�-w� ���BV��lm8���NX{�Ŝ�`�� Do鍕X`��|Y n݁�x�X�����ΌC���
�[N7��k�Y�#��s�>�\jc��BGa�O��Lp�`>,}G|�\����%�������Nz=(q
mbL*��HwUyEg�eȨP�ܴyՙ3��S����p��r�T\�3���U<�u� ڪN��܏�~n���C��KQ��go��v�~*�0������;ׁ�\�/���RY~?ZL,��Q�?� ͢�'rN�/Nm���I\�c�z53��]��r�d�se�rN/��0+��X���y&5&=�0*�\���<3�q�P��q�I(ᴉ	J9*�rg� #�y0�6�Mo������`����*^z���}M��Y$���,�� ����g���o!�zȃx����،��D���B����:����#>��%��G���U�9�0�b(5�Aܨ�1.Nnk(	�ٛ�~���=�8��80�������ꦊ���
�r�C<����%RJ�2[�@�%���`N��Vs����f��s^%���UB>;Ӣ&���O��[���FD~IkX�A�_J٤u�p���$��	e,!_;����[���>�-��B�<�����c�W�a���F�<zK%ŗ�˥�S4�H��>��K�����(�J�䍐g��QEL�ڷx�f1�;�I�W+��ݙ����y�d��&73�H��.��pQÅ�X�S�YE�.پ8�L�������>N�t���ΰ-�.:���D�1�f��5�c�����f�]M��������՞3�#���Yg
.�{]�I�	�b�rl�M����.�|q+��l��ڹ_�(���γ���Q&�� �H��stj�����aW�!��V��5c{��X�>OJP���&R�Ɵx�~�o���E5tz6�����0|�2K"�k�ڽ>�9�d��+�⸾��7ݶѵF���xβ��~��]u�j�O��L+�P)�)�G����e�k�͖'&-��Kj",�,��ڈ�����9�=c0L��V6� V\:��g���ފ�e�*�fE���dm��� �����}b1��s�b�+��ʡ:�9�Ǜ�� �76�ۙrS)��݀wI[�����)�`�f�����H)�z'�л�gG��>��("����P�J������{g��c�}P�6�j�)Ѭ����a��$�F;qq�,�Ux�4M�Ik����������x?���Q=c��B����7!�/�M��0�ň�Op�3��5��j�iڸo{i��K(��p�e?U�I�C,�&5�>Vi�8�D�X]-V�ୠ��4�KVƓ���f+.�q�B�&=8hA�r͌
���;-8�$C�wbz�`�{ĹY�-o���*�E%�g� �̔T�y6���9��5XӺB�Y%z�_�޸?��W��-i�����т���9��ae�"��:ˉ��^���J�̠f�2�5/�(��wB�9���n�RԏZ�U�����𩤼M� ���z��
ٛ	HV��z�t�f0�qM��X�B���<�8��f�;	������[�<M�k����'�ˇ1����Zv9�������8��\�����6аXjŁ�Ru�&s��&���I���/���*,��0<5�e�"QY`��+�(��iB��� �'���Z����%5~ڌ�|mlm%��|D}�$�sFԄ>3���'�|�,с��~��;(;=�Cj��D,��u>^�a�T���Y��VA
�M0(|ǌ�gnܸȧ_��2�O!A,���3�E�I�^���,�(��ȹ� ���| ��^��9"sxx�.���b�A
��"iu��z[uU��̝ؽ����`���Z�a�6"��;��oM����$�mv\T��[[��z%默����8/��2��<���~$z�7���~
�H�䱢Lr�Ӽ�Gg_�=�Ek�3�(ث�l')(��UC���묣�,�׬�L�Ku�g���xeD����1Dl��0�8������h۩�E7�67�k/��S9v���!�"���L�->�I�ڇ~*�/��$�?���N���MH��+����C�d�Z*��CƊsUZu�����n_U�k�&�	j�*0�(�_�҆�*T�juY�ï������u��;�n`H���2�?	�O���Na�������ilk�U��V��_�^
M�[T�d�>6�˯ު�𸩲�"
�܆�E���.���l�u�-��z�1�X��J,7�=�yw�h��g��ť�T�d~�^�y:6BT�n�'c�dX��������5 P�����M�Ok_���=~={��(�1(
H����!�M翗��"��
�"�$XW�lrt��=z�<�N��%LÈ;���3��{q�:rR�<�R�S8A^3��M�Fk�Cf���G��t3�X{��7__�n��u �nuXQEC<&_d�������bx���*�<��֎�ϻ=�M;�W�ښ}Җ^�cX9�h/	|t�'�+F�?8p��yp�w�f��1x6������6��Aq�d�W���Uq>},������e�y���+�o���ލ)͓��?��z�Wt��Z`LZP<�a���òG�Sr��n�O���r��]'��{-A�J��?��Kڮ7�r�L���c/���{���&���h��D�ؤ��zĢYb�9������ჟi2��բ��ٷ��_t�F�:�@���F��IW�@j��~q��B��=o�Ǒ^ލ
��;d�w����7�������Y �l��iu�ξ��R �:�L�3�_�FS�]��`FV�%��6�!�=9��y�t�R �s��1���"1�,"-��N+�W꨼@��g�Y���ךԭQ�#�7�C�I�U���k��2<��r�O~|�e��ϲ�g�M�[�@�z��Sd���8��e�0��}��?h���8�=�(c��GA`2���ȴutUa>wNھ�w��g��WY2���w�^)��[�6�f�s��cS����.�����z���[�L����bt�a�Y�F���AYL!�H��T�p�P_6?M��))D�.'Y�X6�th��ߤ��d��K+r>WxVP�?����t$q>+�էaV�:�xk{��InR�~zj�]9�t��]��Wn���S�U�T� >%��oYt��*6Wwi�iU����˭MJ��}k��a�g`���J*C[��J�̢�K�g&
�4�K"�J��A_ES����6�t�J?0�M�\WtB��N٤%���k��v��jC�:7u �:�	�@�F�Dm8t��w�e�j#��V!�w����zl�<�z�l�T�x���w%i���^�t����kX�^�&̌��MS��W����y�U�ղN�^M�����#���m�V�= �ƕ�aՠ�ySj�����/\`ʆ(k��2�C����\�;��u�t�#(-�Ax��ۜ��
e���,���YI0�Q>?�d�ߵH� "P��\��W�AN�	����?��<�1�`�����������B��Rp���T:̕)H@�A�mM5����#� ��0��=[�:��q.ˠ�.�a�ǹ�E0K�a��	/��9�� #�mڮ��~v�k�bm��JS���r�#u#'(�>�b��l%��8����=�;)�G6��Dhz�jMc�j7c�79 �CuģG�3�5m���Ԩ6GFR<J��(���ZCD�<�10��-�hޫms�l�h7"&F*���d,y1�;�j����J��dR�NG��uV�RS�&Q|�,!�����t/��Cj�L-	�;�v歂�[-�f� ��&t)���ZM%�r�!f������t����Ǫ�4����;;�%+�C[��f�<e�[�e�7=�Ɩ�!��<+1O�����
���7C�<5��9	�J��D>�=� D0��1B"�n��^�U����oLF[�[K����D ~T�
��d�����{֦�E����[R[sE��Я}���D���^D��π��䆥���@�̋i����O�hN
v*���q��U���$��_8�hWq�1/��jV	W��n9y��,!߶�aG�����;���=�5��>�+Ckn�r��'�h��pR	y��T�24}��B�=EQ�`#EI[Ք>�X���Y�� 烈���F7OX���n#���� mv�{�0�l�������҈T9ob}��"}k�U������1��D?���H��)υ�_�~%�oqˀ,��AQ�XԀ�����=��z�s���W!n�R�+>n˽��P�yJ�����xR�Nn�rd�Q�S)���	fך�yxo�e?0�ϑ�^���J.܀�����B��ߵ@|��n�X�*������XH�,wR��W7Ep-�R��h����2�QE.�a����ٷ�����3xS� ~��nE���Zb�#~�}d����3�Ӟ��
���m3�z���7�5�D�2�Hq0x&�NW����=;zO<g����aѻ��s5H0�>��ZY���,�<�K��"��XY��<�g�^bCzR����a��5�@��M�2X�B>1����x�+�#�h5�\�u8}!�P�@��'�!��@�RE ���|��
l�f
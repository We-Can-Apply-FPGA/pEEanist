��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��ɳ��a�i�������L÷��������Fͱ�y�.��+2{��,zf����{�P�=
��^.�
Gsܻ����h�N����l��!Ѵh�����d�u�t�!9/�f�=b�:O����}q#�����ʎpH\Ju���#y9?� �y}��8�6<b�5-�l���Y)|A8��'��|sx�����g� �
�N� ٺ�R���L��0��eHXׅE�M��7��o�hMj|O{�	���{{C�J���L˂8D'�Ʌ����%t��z?k�.�l�]�'�'^���_ч��w�(���[g�+���V��6)�gc*�^�`<]w���M���7!���rZF�^U�"f��ď�
d� �l���V
�uS�;���n6�h �S����P�}3{$�=��}�������:��KX�23(��ӎdMm:.JN�����|��pF��$ sdlI �ԭ=7�X�{*C@*��jǒ���(	�J�ưS �<�F�G�O�{��gD[��g�M��B仧\K�.W6@�c��yÀ+��Yo+zJ+�6A�-h˪�����vdA��\cu�e �a�RfAW��?D��^�!v��sP�f?	d��n�Oh���5�� ��h�¶�Iǣ� .�7=��K\���\<��dG>޳w%�9��S*��뻶����6H^�TH���|�+x�#�n5�� ��-�V�����Q��`���F2Pe�0��y�Ot{g���R�'�7��"�tP�{]�Ǧ�="l�΁i���,�������������6r��v��|��G,��%�er��/g��k`�5J�_a1P1��T�Y�[5��}�1�)��\U�Q�tg|"k�o3#��-R0�1���(7e@���D�5�b��9nQ.ĎS�o�yE}�A�Bd薗n�b	eNR`�Tk'��z��C�若uj�&��d<b"s�a:lǤ+��:I�H7�K8)�z�fH~�{,:�˰>�E�qssPlze�3�ao�K�3�V`���Y08��]�)Pc�ȋ]�C�h�(Vv#�!��H7t#�|�<}0�j�Z�����R��]��}7�fhӓ�V�(��2Ή](�L=��7o��-2�\��/Fk_8_Ԩ]���k�,-��>W���	Q�jt�h��O�>��tȜS7��e7`���T+���s��nu��޽FT˔�� ��)���]�����"����LhԵ�A�j�fϲ�=-	Woñ�TȄ�C�<u�_'RƄ�����I��J<SC�A�[_o�"N�q�����%�f��܃�����)��:Z�4��nK>y���Y���9�+�E��Ȑ�>�;��E�]W��Un��Y<f= ^/9dt�w�@��J��P�P7$<O>�ޢ�yER2��YX�+]U�}� �@!�o�p#�U5��"�%��4#�|��ȵ#�r������"rS�N�BY�r�Ri+Ć�H�  �d�b��m�%j�?ۥ��e�-r�,����:��F����
���s�v�2�LX�< K����a����� L`_�[�co�����R�1�����<�	���Z��\�tYVm�kP���w��oé�h�X�`\�fҠ���+1恣�E�5�H��:\�>�Դ������0J��J�����@�
���������F��U��sM��'�o�R� ��Ɯ��a��{�|ت��p��U	h��[�w<3��)b��I1��72�9h��u�?qvB�8���jB�+���.͋i��垿c�Bc������z�*�&Kӽc��t֡��a�HT��D��-?_�V�&X)$�c}��ٹ��m��Kq�[��;�jw��؜����V��� Hxt-�}y�I���Rtu�Y����XӚʹ�H��`����R���s�o&��*u��D�~��
k[H��VGZ��צ$��@L��5ǈ24pU��/iilz��R/�+�&��j��Ao �	�	I������ã�'Bo��摐?}>�
bT��$�[ɲ�������5�ؚh��V��+Po��	@!��N��\�s��p��M�Q�h������޽��A�n7��˰dZ���.K�U�nZ�V�-F��#'QqBg�`�%x���L+n�_�D�BF��`<�� ю;>e�����䥱�۟[�?KQ�{q��??N��n�}�M6P~�����R<%��{)��v�^���~t�@\��?+\ �eH�li�YB24 �2��D(���Z8|h{�"�{�rz�0]}� h�`���v��{��H��Ap�3�.
�n�FO�_�40��@��rr��O���'�h��M������Q� C{���ӄ�92Έ��WN�`e��
YO3�b��	�,P��ߒS#v~�f�|����a	�|�/�M�b]$�F����E��q���%����R�vl̋{�#�J���|�>�#��"�]5T��`O��{�bp �\�v ظ��h'�?Lm����n�LS���n�iivi�
Y&w����
1.Sx�:ڢ�dڙ���p=j������}d�ީj�����t��橛}A�A>n��1�S.��6̸�F��]{����-exjMGNb� {��M���S;m�ݦ��{�H�l��Ӊ95�B�Z檈�]h��fq�D,�渉��n�^`yHT*J���^��x�c��G�)�E_�E�UgJ����!S�� 
�I˳�O���_�a�ˠ��K>�=�Z�$_���\���\la��0$�VB ��-�9ul�2i�u8��J�ްyj:š����u�Hu�p��b��E��օ5jf�r���LX`���Vk;~#`'�F�U�7ַ�k�zXJR�:ĳ��v�h��W�A�rݥQ��C�X,���9/�rgБ;.a$�p}A�G�$�_~@<��ka�=H��@ ��V=�U�(���j��
��u��Mv	�'�M���/�d�Դ�� �-�K~��������`��'S��Ի��,��F�#���&�y�>N���6�D���k�_�����m2��Mi�l<�������s��RO	{N���
ɉ����G&�8�D����./�u3j��]�n����+̀�(c��5���*3�:��t���+�rw���-��s�:2&J�9��iC����g^*|X�)d��_��Gᢒ�������d�	J��;��G�������]֑�2���A,��%R�+���������jp�&�/�L|�9b-0���#�P�"��c��S��Ai.s�	�J�l@Ԇ�F��K�Q�!P�ux�պ��G�������ͬƟA�f�$,TI�[����g�z�}��)�pٹ|Ep��� &>?�U�>�)�Y����?���4���sK����Y*�\��-F�1Y;�?��@G�Nk04��Y��xJS�1�W�f�!���ݱ/���A�C�WGΰA�杓xd��1$��2���)R�x%��i��D���-#t���}3�M) 3�D���T�p99�,Y��'k�."/b�:Z�}~�O��tjO����|t9������imj����|�m�l��_���q-�^'���J�<��iM�[h��@�S����B?��y��f�<	�Ki�m@,��6�[��	��U�����%�D��Y+r�=�Ζ6�v�v��H��c�� �Z8��Q�8��k����p��ؤ� �u��or��tS3P#-��_����\)CX����jxޒ+j���H`'v��i�!��kD!�;-U[Z�N,M"���`K�ia��Kz��d�)/_$ųW3F����Ū-�W��~����L����-$��p-m�{�O+�o?���EY؁LT����b��v%�R���UBs�&��(-��<f*㨟&,�.5J��c٣�W���ђk�Zqvsٝy5�+�w/����<��7䠮�(�Lt.�
ݚ��H��,R�b��,� �,6�:�����v=��ֆ=�p ]5��s�s��i�e�+�e��,B"��W�Q�D�c2��`�Q��Ѡ����̡�`����tyLs�b7�3uS�Bw�95�F��GHP��Uȅ'0	̳���d�@����~4���d5��0־ʱ8ሦ�-D���
����,�^�8s��yBq����a� A��\��0K}� ��'��	��y���7I��A�}�'�4TG������M\c�7���3?>M=����&��ʫ����?�q������"Q��~����YU@�;WDX2�a���>Y�p���$�cRS�39��~GXx�'/��f��L�%��34��/"r��k>�i@�͟�Wˏ�����/71�P$�b�Y��r�r0!�d2�����]6�>��Z��#�>>��	7��p��'�<�Wf_&te�,V)< �(�Zc��Dg�49r�KkX������˙�o�����|�+j�W>��'�ؑ��T�@L��_��O�K��2sg���(�۬���,�W��G:�_T�G�j�j��a#�q��G#>颖��$D(n����:��G����>�F?�t[ɴ�R��l�ަ?'^��C�:ɤg�F;�$��	Q ��E_��O�#�V�JT}���J�A�g#� �QD��g��J���o�����C�;-|{@U�d'`��|�j�iH�����4O�Q}�ȸt:{.�T�8jWI�@1��zz��x
�e�����î��,B�J��0	�`5��*3�7d�De��x5���V�L��1+�eВ]���N��-'\�'󤋹5�'��P��������h��j�$�=���n8��{�w����ԡ����/ͽ�������|�<bpk5Q'<+��}�w=M�"��/J��Kh��i��fvMF�u8{�_�<_�Tf����&���<6�Yf�ٸm5����������(m���d(K�F�_2Ym�Xlp6_5ؿ+.���^���Q&DC�L�lb27��1;ށK3H]�<��b��1X�7ה�\���nU��7+��<U�Xwҏ���
#�� �q2���j�kxr���#+2�:��^�˻�.
v}��Wc�]���eĦ��6��B�H���Sw������g��?q_J���W�b!k'h�> E���]CIp�ƩvE;ɥw��L�Y\�)� �
(��2P���f���U��fy���6�ņ��&/�][���zo p�Oa:V�>h�f���|/ A6A�a%�{
��F�rOK���Wf:]�Vj	L�ͬg�ޱ/>���9D؛���/���ƫB&��*�|�� P��!�?V\�h�syZ+S@���¦��K��I�y'�G����_AU�VH��9)"��/j�ʇ0�EH[�k�l�y)�
��+�OW̔�\�|�ز/OrQ��va�IO�`cf}��n�p�*�:��[�X�_�SJ�?۬�`C������Z�+NDh7��i��'�$�`JgV�v/R��;���`^��s���"���z]J����9�ޗm�G�_�����fN~棱x����&}:�;���y���Ͻ������⨋���y�b�1��Ӄ�?��)	�7�=��:e���)�b��Gl�kw�ˁ���6JA�3i������l#��h[S�M�c�|��=�d6�"F�;�%�VpS?i������i��V8RH����`��P�CA�Mu�.�ˡ1�}��!k�5�kK�?z�T�4�n�{=�ZLy߻�x`�/�7�_��5��W�4r	}���*U`I�w��9�D~j��2���̅��^�i�
�B�]�A�E}[W?;[~��6��|ɨFA�p���Js�{N�ߚV���H�����3�l篿��xR������&Y��b��~�F���d{��n�/�h3���x�F�y���0*4脺PCEPLC�mG��{�>g/�A�R�Ռ8#�uڞ��Q]��Y�9�J�pQ���.֒�Â'�u���ƈ���¨����U�By���
��c�J>NW���"�^�7� 
a?��31h��N�z�i�h� 91/���$;0��QP1�D	��&Z+�Ǌ0�R�/���z��ktjg��`��p�F����hՏ�T�0�W:a�C1�R~FU�.!o���P=��;�5`m�9OV��)7���K�\��]=b�����v[ unBʺ���@�	[[������X0?M����
���-AM��ͩ�B�2Xd$�g=ܰe=^X2xy������sV��Ě�=�"��o�⯛�Z�dԢt�=�6H^Q.��`������eu�F>Q���Nr���@��H�1����J�Wz#����
}"]S�K��3��lV�ڃ�a�`#�H	���1���V��R���	ۘb<�,vK�b�0����j��uK��y��a7IV�=����:��ޱ؄&�o���J<�,t4Е���ۅͬ��u�ơ�iXɢ��g�Kr77�j۸�8��CM���㛏�BGu���솠ַ8L��\,��+��_����L�/�4���3��]�ƣ����%�ͩ�g�O���ѵ�h%�����ƔO�7D;�AB	��@���_���`�,��*�x�A��#Tֳ/ܒ�z'�ҽ�s���0j��N�F���K)�"�����~$���Mx� ,�L�mY�9����z�l���K�	!��5�X����	��3O��}h�������SzuG S�qJჱa��V�p|:Դ9J��#�|��o9VA:&ocw.�G��*w.Gj��^J����u��IB#{T>󬲼�)�/,�i��Q�X�%~��;�/56 �2%'.�)��ՇW��?u=��_u�|�m��0�٪��R�W�kϭɽ7;��Θ���B=kw�\�(Y�"\��E͘�,Q~JdbL��[�p�Z��q��X���c� ]��ێҨɊ�_h����3��$=�Z}�H�%>ŵ�:�5��2]E̓/n�30�"���'Xu��]mO��Xu�������[�HK{��h���*N�&��0�6��K?�+d�-����d�7��CS;�g �%���+t(��~�O��� T�I_�0v�-Cπ�im����+��]��S�(�>0oz���"�LU�F\�B/L/��O2:5)j:����|������:I�;M׳Dvl}�\��� ���Z�Q��v��8�K����*ԉ���-)�b���g�;|d�tmgőșU������ѵ�����42b�_|���
��Ǣ,�8�(�W�x��;��	|��6-���@P�/����qW���� o$�	�aw��@50��M/��V�k���i4�غ%�5gVk�\�RMP�r3*M*)��7�+�lq��a�8n�~2��V�B�c�Y�b����A���ﾝ?��#���UYi����d r��w�j��e�Ld������]�/�4蝶�m�[�3�-ӑ6x	��-i���J}���;�`� ��5���/��S)spq(�I6\ܘW�)�u�B�~�9�C � �;	�9�F]d��>񽊰��Jͻ��'�[r^«\��f�BYi����I+Utaqia΃�zƎj2��а�J�{��Y��'x Z����ƜNf�rPm��<�Yg�h�/��ZNT�۸f�Ds�*����K����vz�3��A3����q�0�9Y��Gt���S_���&�d����>�;�l�B8�>t6�����~�~�i�_:�0佔.<�����\'��K]1����]���M�_º?���SCd�X"�Sn*Ɔ1��
* FA0g�c�c.Q���[Bگ�Y�-?e�;9���E4k�ɟ����s�l3o�� �1��|{_�(��h��y�Z�8�k��P������є���`v1���7?��_�G�,J��UMB�_�O!�w��2�Wcya���z���IS�b�N�\W�6B��|�r���fX���]^��?G���@�M�k���y�ˢ�1��C^1�?����Z�s��5b}ߦ���xH���u��b�Eڜ�����/���xw)�?6J��x�.ԅwx����8Z�΅s�́�?�P�9�Y����?	gDl݆I����Q]Q��֞����ȱ�բ8$�@#(!j�T���I~b�oN�^�(C>�g-	t���)�g�=�&��N�1�V�=�k{N�?�E���2�X#����k�X��{m�
��v�f>aE��Ƌ�U���i�P�p>���0���ڇ��fS��Hc_L ���3�l��Ǧ\��oiǺ��`����A�SJ��oM��\]�<s����?H��^��Ft�q���
N CB����	?U�T���qb��*X�H3{����^I�p?��\3e���
��;�����6��;1�=��at ;���F�N[D��P�������	<�V���Ӗ�m�i#�A�ff1Mz��E�6Ѝ�j2��
�2����@�y��#�9=W�'�T?q��wijM`d�kW�3�����۝p�<ӧ�h��h��8Nf�[(���$}�[[�6id����1xC�V?��7�c2�K���nV���6s#�����M�z�k�C�K������r$گ�7��w��zP�������!�P�=��S��}PS���{x�>��Js�^�̂rXl��t�>2��|!�dr\+�0��΁N�F2I��ץI�,'�O\�q����Z�)��e��T&��14>xE��c�Ӧ����p1T[� }+����7�����C�3���8Nn�S^�YSu"_�E�d�@9�Vι�Tg�Th�n����Mw�G���'�d�z������h>Vݜsy��������Rw�:)
��m�g����@��p疻�9ݬ{N��my͐I$���E���"�3���!hm�1�K��k�
����8��c ���¶�8R�){���Ʌ����M�BgC��
�z���M�x4�M�Ct`c�k���)?mP38�p^+��h�g����){(Q]�
�����izZ�����>�R0��8����ˍ:��p��,u�ܒ1cP�����b���}x��>�3����b3@���P���b6@�,�I2)"�5qO����L��rR��T�,+�[�[��~�B%e�7���(�т�I����E�v�� �H�8�$��s�p�4|�M�OQ�Ŝ��%wX����X��ƭ�ぴ�^���V(
�Y� ��!OL4�7�*.F<H�fד���8�o-D��}v��g��h���hX���I�FC�z#gf�l�&���K��}ϵ��	��^����+���;���p �N�CI\{͸,ݘ�ͼ�- ����%St�����v��� ���p~�IN귗�C�j��Lh���}���2���>%(�&ֆ��tn�3�UO��g��ųN�K�x��n����,�2�@rB�����=�ysS=^t��VN=st�标�N��9s$?B~%���g�*�F���Qc��)]�0�6�D1�H +k}�ՠS��4B�� \�iS@ܚ�p <�%(v}���.�dX�[0�W���,�JE�*v�/,	\�teO1>�� ��4���8���ԉ���	�C��c��£�߳���%R����甎GrhJop��em�sXPt~3g�*&��	��k�_��Et���`3���yA4p��k�I$
��kvZ�.~ ���G��v�䪇C��xn��E Xp�!u�qP�4R/�Nߗ6����8G��Nr�:�,3:` !�M�;n�,�.W.|��?����l��(����)n��u�n=.[;uűVD���H�ѧ����G�H�F��=K�T��O��GAa���{��9�oڱ�DI�A��v���,��:V(m��T���|m�˝��2�4�x��p,,���C�gY&���H5���6ؿ�(r(�<j�P.E�d�~Y��X����)��8�w.q�f]N>�wĉhDp�;�LX��v��vi����Ø�&.d��9�7'��?��xUF�\� ��D^d����|H`T��5�e�ȩ�l]r�<�%�'E�v/��_�������1p*L����cYΩKW���D?C�����X�Թ�&�e=&� o�B��#c�X_ x����X9$7.��>���s.[�W#����;C=�2/v\� ��N�eJ���p�)�W��Z�g^N�d�F@�w�����\��Ox?	e��]���T�"�|2���PgZ�����k�E//�vX�u�%\�Q��:|O�EȚ��lu72c[Bn���$
�f���N9�秏A9|���#����� ��8�b}�����g��8�9���hu5�i��(ܡ�R���.ië�7�W���y�v0��z��6��9w�]�;z%�R��=%as�}Q&0��P� ������#�+b�v�u��R��e���Փ�>�
�cK?�+ �|�
V2��(���jO�3�_�F��Y�X'��G��P�O��e���%M��U|H^cT�}��'a�K�aw����b��_( �B�M���D�w6���F�1лI<;�n�q;|:��1L��*����Hr�s�77�� uQ�V=����:�o�ѥ ���L�;�I�5�dR�Y1_�&��~� �1�3�j���4�W+䞻�_Ri�B� `2�N�$�(3�d���u���wR잞�h�Fנ�����6I�.�����`$ں��������j����1����de��Lף9$�M�N=��(|�L)����PȬ�Wd�ڏ�{�Q����2W�(:lKt��L;:1E�%$��ꕅ<u�nW������b����M��:�7�C�q����������i��q���ڡ��V�?����Il7�V�\��%��%'�.���!�s�eh�a|�ϡ^��<e�wI�\3˥i���.ˢ�Du�-�η�SR��jsDB�&%�I�5�	^�C�C65(Q�Ӆ]+Y���k���d�i
��;:��� �XR*t:�#��8%o, mt�Ck�$J�
�?�\=K�J*���e�+���O��P�����[ӓqF���lG���!��Bg�'���B�d2g`9ѻr�!���6%�n�M+��B_j�p4�)+��ОF/ u���s���R�d/��nU�y�@F�.�4}����T����q?�Nv)7"l���Z�����=�Bh~�.wDd���|��(�C�DPd`���S׺Tu����4D�`�皖J4L�儍�%��.������қT9�\l[�o����"�P���������Q�%�F͡�C�9�I� �zHa�S
��>����E*���j�_v�������rRF�t����Y>%Ҁ�+�����s�-�3����Bk��֜�TY�Y�j��i$tGu{�+�/�c�>��ۼwږA
�D���w�>|�|���th�㪤G�̿9EF�N�xE]�B�C�ݷ$M��;ɶ�^:T���w���q�|�mvd ��q�����J�Z��._�#C$ܤ=-Vգ�
�j2hO���9~2C�cP����q���8�q}C`�}��ڮ%�r~.'_w�K��6	��&��l�_��b㯛]m��M?N�?`�LͥY\��k�,΁���h���˰�zx\[A��D���:���#$�v+�7"$o�8����g?B ��w���!ƾXK�%d{�OO�By���q]��&��eί���ePm���=3I�ty�Zq�J�|<��ڪS$×�yg��gl&���<���SG�/�A�}m:̌ش����n�n�ᵽW
�\97��E��X�T#�FU:Z�H�'a�����pj]Z�	��V��Drwb�9�ԉY<Z�hR1�W>Ӭ��]J���v�Tʨ�`6��rZ/���Â%�{Ej1[&��� cww"��0�>�������"C#*�e��2�Z�dr������<�t����畠!'�Fm�%.�%B)t���E���Qï�c���!��j���>j�$�~=8��BzC�v�s��G�{͆� �?�B.#��P��l���Zub�.�e����WDg>0�X$1Y~�&6��~�o��c4��*2�6uh̭�5)�5�b�l��$�TKo(��vXB�O�@�[j��\u��\B��zv����}�0�j�j���<���ѻ�Zas'��F��p_���#���uk욺^бY�4���wp�\�)+&������7F�q�Ҏ�C��\�o�9\��b�*jfm��?Y�]�d.\⽯�����������s�m����ʿ�p���a�>vW��	�O��QK0����C��IF{���cA���o��]Y��~� �!+�s2���'�'xfN��I��sk=M����<�nĿ+��0"�"((�v��\1;�w��Xv�k Wn=�o��ZA����6��I�EwM�/�qB0~n�4��m��LB
S8��;q�o}�����nc!ַ�p��t�F[jV�#c����}�e��P�h��#ӱ���bW,���ʵ�_G�r����ۀS���z�0��*��.�1`��e��H;�
�L�7��'�@_��M���K��L�2l桠�w��a��Ul�Vo��NtU1�W̕��[�΢]���)�7���rm�aaI�ʪgK�X��z����-
��fU���4f������2N��Q��ea���5�BS9�>�kS�,��=�n��~��gѸg񣔕�n����-ON�2��V��C((ѱ{�0�R�' e�t���j��4��t����@=ў�ed��X2=dzsj��W�MkSo(�#��=�ӊ���WdJ=�{40��N��XF��O�
�-��s��A)/����(��3�J,U��Ǒ�����U�����̢�6r��e��ٲ��vA<�̀���|	�s�ʈE��#!/��u�p��8F��lL,L�pF����������n /	 m-�s;������[�Z��L���6�3���x�~�@&<Va���&�z����2�s���3L���<M����,�u��#�e��!�o՜���N������ҋ8��IJo����(�C�H��K3�g�
����	5�_̇�F���"TrOgi�  �o�(��޽y�^@�`�թ�k���x�b��Ő�y�V��������aq	)Qz����j�!���?h����\u�.5��{�'��0�0���4�n���oe�j����ṻ� �"��(-�U��AI&Xd�t�)�͇�4 �k�J�l�]q����c��k+M��p45����`�fĕ4�c )5�<���b|�0m)g���u�ryQ�Y�yE�a�) ���0�È�x�<4���7U���Ax��n9+ˎz�~9�Wm��
���֘&sqm����H�:�n&�'�6ٹ�'w�o����%�Es}tU�p�G��僊\��A-���x=x�6..�!�����L����::�\�El�:]����R���Ov�l��GE�J�;Cd��m�Pj���x��
E��<���Y�r���'ǯ�j�6k$�y��&�.y��i6DP�ϑQ'>��ed]�΄������"��4�d� i�e8^{x�Hu�V�ۃ)�� E���#���?y�����/H@�2Z�f�Z�4����!͛����WB����L��[gcL���T�~Q��Fnzrc7�,gAb��4E��쟸b�̥��;�{(Ζ�}<���31�`^�C�!:�i��0�]�|��5
.ST���gj.P�h��m��#1\��8����K�.��{��%ס��ɹq�:d�W�*�����^q�} �?Ó�p�>(ߦ�X��@5~�~L.Q����6˱�&�=A�E�|:'���5���~�i�pRv���'��2=�>�]0��^oJt������@�̎�i�{FHA켭�F��Z�����%�&��S���4�>:O?�~]Rv^��K��7:FK4�}WZ�d)�֚J���q�$*�8v�n�=ъ�᳔[/L�ޤ��5�5{��A g
����~�
H0X�>���Ѝ��Ekͷc*eyO���鐧����1�i���G��Յ7}�"���?^��+�t�ԬM�ȅ��]�s�$X��1���P/kEI�C\���&�X�S��у��U�u�yȗ��,ޟ��-5�7 4�Y]}��NE��5b�F+�0al�#F�1���\p��$7�D��a�wqp�T�e趌�_��,M#$���ϫ���c�����A��|!P�j��æ�Xtc_����⤷0uu�θ��>K�Z+T�0�C�7�E)��e������]���r�qP�R��,�Cc��JFVՙ�Q=\�;�y�U3��:��ȕlƗܻ+�r�w����Ջ�<���Ƞ�Y��z)�P����i�ˢ���Lf�'	"O��	���|�����}�}������ �t;�F2�(�gx9������s9����]oc�Į����M3���^Q���C~K��F'��wNG�`~���s��~�Hw�?t�'$�x�{��b��4�&���Q;,^��`�`ҩ�:}6ܱ֬���$V�=5���"��A��U�|щ�#j�L'sN�ǰם�����.E���)&
~)��(5���^rԒ}��� I}�oa�3��D�rOQ_��8M-��IQh8�G������N#�K�"���neY�S7=�@q�h��?��8QR�]_#�h�����kj��
��\�^
�\$�&�VGL|��s���۝@�IپWh�J�ն�6� ���=J�s�@��"n�7{�`��e|�ۥ��'��¤�ɟ����B�϶�����(
"[k��ن���R��~�0����!WW�ge���b���T
�q_�e)ٲ��M�	���na��Ge�3���^���idKt�u�h���S�Q�s ��,O?!Q���`@�u8\����
�
�M-+g�n�w��?`����Rb���X>�y)arV�T�Eof���P���M㸽v��AH,��W����h'��yEe����~��s��~�imͿ�o9.��Ĩ�m/I�|]��s\b�T �;����b��y��9K���Ų���؟`1
%���MD�:~�������I&j��������(]�i>摾b��s�O�y���C�w�(���\AM��h�q� "
���cmѳǟ��p��˾V�h�`w�� f��`�?֋���վp��ݰW��k�N��Ma�L֗�2��D郼[�:�pS�����0:�j]��#��^R~9�(͒Q�i5����YW%yۄ��������o�!����=N���!��\T������e��~FK5�ew'Y���t���A?���;>����OƜr����s�٥	�P��	��k8�U����l�h���t�pUk������<(�yİ�q���Y`��_qͅImկ���MU�Z?���"y"�H�ȎOH@���D����tt�:]��	:UbVI5��mt��.��F��7�;G�M8����h�;4m�Z�1�^�Ƃ\	��*���|��NO8��޼��z�zl��u!�o��	0[�Kd��� ()���+ǔ�"/P�g�8����h�ȇ9�MЧ�Yy.�&��_��G$�n�M�]��z�ɏM���7S��s�F�����@L"�%�H}��iq��Wۜ��<ZB��Oٔ�J��R����
]�uht7s�t�7���P`�������� �p��;��?y�C�H8�}��{��S������9w�4�g���h��}���w�9BɘTV6��"��J��B*�Lm�ExKq\#CC��m~ӪKŞthC}�{c�H�%�=:����N4�D��e	}L�-�%-�S���x�|�Su����K�)��_��~61�T��������pk��<WE�V�s�JM��̎��˰��6W:(�W��˕i���\`6�Ѝ�S�sgO���̻��+{��W���Ł;9C�^KB漬��b$+��f�!R�[����$��e+S��!V�� �����J���.�t<����M,@-���6�.��D�p2(^����������͓ϋ�����s|>j��⢐O���ƫ���k��#wq��:��@d@l�ͪ��(�@�s2n����B��ԮC��~\k�fv�Y~IJ7g���vݷټ=2���g��u��>�͑Y����ϽB_�����-<�^�a]�g�p�k����Q�$����g颬��]<��ON����%P�}�1�� 
�Ow�(�2��Z^�a�������s��a�Fl��r�h���� Y�ʕ|\����ԛ���&�%�1U���#�����m�}=��C�[�:�w�f��i���A�̈�rQ�{�<*��*w�p�W{���b��I���=G���jsF��փ�Z 휊dg�b`������4�:z�U���"��|�)���Q%n�Z��JI�N�hd��r]v�R��9V+*R�Rg��r��ٿȳʪ��C��*Y��F (
�h�$_c�V���L�,�8�*���F�a��p�/@U\eN)�aߏ��U��Q�1��G���~���}��u*G�i	���n��ȫA[����!�j)���� ~3+N��r#��2p�:�ƚ� $,T��a����-��ʝ��͐�W%0Õ�5��Hj�7��* �6o<d��E9ry��IoA�->�����kfWIC ذWj��cQć�
���Em���w.��+Sr�Tf�r��#i=�P���Ӿ�H�"dڃ�c��p�/X��{�TPi`)a��M[�@��I��5y�<��pj�+�C0ͽ��$^AÀ�_���Y�+�JP�LT�
Z��RKآ�B�+���@�וr�x*���E�'>uL:]G����^V�s��\���"�Ԥ�**M�`-3�"��kU�4����A���m�v��]��{�E�KB}G�=VXV�T^��C��:�{s�+IP�8r'ȡ�o��1O�"f͟=�+<v@%�P#�V�/ X ���ziO�Ǝ�q����s�e��4P
��ِ�WM���d@�:�XUs��G��`�M]�-�0s��PL޷s��%��k+�ɔ�^�H+���s^�o���:;ߕ�E.�*�!IΆ�/�LJ�����b�~ԝ˙������Np����_��ޝ�_��8<����5R�>{�)����I95 �,Ғ�C,_�WDP���	���Bi )�5"�����f�]�����/ �{�˃�Ƽ#=1$��bi�N�������~�wS�&�����ωjL��d�
�s�MhB�m~5�moԿ��	W`�{���7����� q9������慑�����f�M����2���A6��A��?��#��Qi�xy�
ᑴ��\�৩�.h����U�g�������u�qé���t�׾lf|/��H��H3I���47�ﳟD4je�'
f͢K��ݫ7&n}���f�]�s�����b� Z�-��f���%d������UI��^w��Ӥ(��+֦U�A���dv^��������N��J�}Ɣ�Y�ĥ� ��(q���am*�Y!�h����,��[�V�'���
w�.es�!�W=f
��\��v�i6CU'U�h���b�E ��ӱUYbG���j9Y3S��A�躾P��?�CRF{��M3��?�5����Y*��5x�#�ުu°�Y9mW=*6��T/����8ėJd
���`�]�xW66A�}�h���Bfp��EB��n��yQ�#�Z���y�"2��� ��˳6�C�=�P~ؘ���
&�h��J�~z$���.�P�X��i2����Qd����p�뗸aX����Y�~E�@�
L�PW�>��Fލ�
i���s+��2uU�E�UL�����1�������O���|޺GDT'�-�� ���G@����>��&����ss֪��4�-��[j�w��V9z8����»�������q�K�S�i�y�u���~���*f�y-���Q�*��~@�@��)��߭g���~����蝼�#���7�S}D ���"x��kE$��M/ ��ѡi�����$���g�u�8�8����%>]�i�|�"�x��f�H,�כ��ޚ���t:������Q�,x}��*����E�u� �;�i�z�Z����>"g����Q�FlWZ~@.<��N�'
��0Ub�9iŲ�|(/�P���u���-��~���AK�.�ƈ�LD�B?ZV0�o���W�)��n`� #D� �]����x,'��t�i�PX���hLd� ��R��Q8������lvCxt�\��{�;Y鋖A��NNJ;� Q@�K��'�t`�d���L.��	[)�r-_	�G���&)�J<�T��z[��-n/��Ʈ�rb�Ŗ���`�c��/��}l�� ��f+8��/�L�#�Z�02F^X5@wINK��4eݿ����漿�hda��W'��J�W����N��5����]�_|�#4ɨ�����qV0�:
o^b"�+7���;�H'=?B�X�զYU�M��`a�{R�y�oD�1��h+M�Ku�~��=L������Ӛv��}�7-=��mu�5�ceN�N�5�j�_%�E�'����!s>��R[>�w_!p�
~O��oaI���q���ƶ�]�]���:Uz]^�� ���X6m�:Fm���;�
csf����{�\o�_�\��e{� k���c����D�vRƅ~��/,��{1tx�A���1X�ԓB��%IP��G���!���OI:k�LlR����?��&!h"	F%���,/$&'��KR�
W���a2ND@�s�b5�D	����M�����*%�-���n�`�	�06�WqY�\ s?`�������~��ҫ����R�A�|t5��)�r���P��W�E��k�h^�Ƃ�<k��<�f�����ѯ�Z j�c)p���q���0������WsI� !��r�Y�ÔMm�na)�OO�|�u[$2r����j�9;��8�v��Զ,]�a ��n�¥�dCO޷��-'T��T>ԛ���ͧ�{	{�r�Jy��X��[�)	aj���7��Uc�2�Bg	��7�x��ټ�:�&쵼ы~TkP�]�Ǝ�y�M&��s��Y�Tw�Sq���_*}6��0�E1���A+v"��ō��>�O �Kzd�8�pjl�D���q�q��'����g�k��(i�����`U�W��[1�E"�Jq1 ��p�a�gǮL�O#l$}��B ��{\�k�Cc��)��������d�`�Hu	xwS&ʤ�eyT�����D�����Ŏ��G�kyOov�g���~��.��Sk>�0�a��Ba�=##�5��
���C��+�=��N�!�\�1
]Hd}����jJ���"�����ٓ�`�U��sbqaiM������7�=���.��s�Mň�2r�d��9���Os�p�:^�������!��
_�|�=t����q�в_ѡ�J��U��n:�5H�Q��-���%��C���}M��~��	7���sJӐ)�����w�J[�c�]�
r�:/e�~�ZN;i�UUrAd����n�נ�;��o�Lj}�:�[FN��4������m��T�+Qe�vX] ����E"� �y���G�
��y󸟭��f�JQ��ku<[3�@dFS|�h��;����U�����KH���ل��X�q�wX(&�N"���P���P������pG���_�|>��4��Qi
�������hbp8�:�M<�U��#� q�4K��\�cѺzn�>�b�=��I��ͻ��U��%fQk�6�&�0�����醷����}����m8��Ə��ō"dSǬ���iC8Q�����:�Qls�eE@P��a]�	���3��9���n.8�[�Ů� _�SrK�F�a��zU9�qSY���?�G"�>+�-M���VpWNe(^F9�b��Z�H�~R=���r��u*�>H��1� �� ��db�턷?�)ʕf.���x��~M�.�F��rT�eҶ���%/����_%I}C���W��\��]Y屚Z�'�+Ϡ9.��t?-��C 5g��=H� ��߬=j����ˍ0�M�O��q��p�����y�_�S�[���O��;_�M̜`@��|��̓����.kQS��Bp��sX*��99<�H� j�����X�K��t;��OIϋ_�E�����]��_R��ĉ�宺��`˞\�<zI�w�r F�xP>-6����q���>���E�,�>�Ee��<���	����I�K���țɩ�]z���?<�g-�����qBE����()�_�4�b} Ϲ��C���NR����;��'Kp>m5=cJ���*?��P��Q���Ih��D&n�6$|yٷ��r'572�Q4�ӪZ*���)Tu������r��{�(�u�ʍY����Χ�߫�%S��>��RO�[W^j �������v�3��3��}��(��,h�uʞZF� q7��-�-�����}��\�]дJ��>ظ���2���%0�������ѝ6`+�}��!nI���+E'���٥�爦��GAa�KB��� �9��R&���-i[v���k�/&�o��$�D���RTW%�/t��5���9f�d�`�Ӏ�۱�z���o��=�Fܗ���Q��wۨ��#:���T�Qa�S+���r�w�PoV�\�JxU�����I�/�#����+o;ʀ���9q���
��
i_n�2	�H6��гz�`$�gx�c���&���u�~Z>K��G����,��,�=Tݣ�)N}��{�@�����DQ����<�a�u|��֜�Gg?�"Pc�g�d��~���]�䃯�b4���A�#,�ɸ�QW�� �$�]Z�����Vm�]��`��"�R�;�o�C���H� z�hr�[[n��׬S`i,+,[I�A�E�70'cd��D�]��۵��˪�i��win��I%�U�5�R���Ȝ��!�S�s�>y1������$�1�aY<Ed�����߂���ަ� ��L�D�M�V���L����K��
�S��cl-#d��l`l��\q���{]Ac�r�y'���PC|u#�m�F��`Q��ϱ���e�Թ�7_+�ϝټ�T����r^U���a�+��F�[ծs���DL<�����آ�L|M�]d���Ӄc!?DIp ��b��L�!J�� ����� N�#�-o����]�R}��������a�	*��u�#��Z�^vo��.�9�md1 ��C�Ȉ��"� �>��_:��U�l��;�XǴ�(׊�E2��d7�	�TA�ףּ�N�p�EI��G��)��[�r���fbH���*��b_���AQ��	�8���`�Xб�����ͻ�y;_�7��f���c~�]<�!���𕂭���g�[��R��#�8,�]�x�����S��V�m�b����'z���kW�CL�
�c�\E
�8����)ܕ@i���a�K�I��|N~,/�LPiU�����Y�u��	�.�R2�@m�0��TLP�`����+m�,rG��$s�4��H��KQ"�4����{�'FLv�Z������F����L{��E|���􀠜;>={�$�)4�L>�̥?=�,��w�	%���d:3)I�ã�!��O�<�#_�5-L�������a�>�>ټ�ӳl�-�#{��m/�� �����;��6{%�� ���l=��	k@*���H�&T�\�f�R����u R�d�G��2_��"�H�4�g�N��.��Bf��
��sS��wG1�0��8���Ƃ~�g�
��V����!�<�^��>x� ?d�q�7��*�2��bT8��}9���ծ���@����E�$�8���]�HB��8��Cs��U�-�,Ǜk��{6n��xR����ڦ�4���	W���:�DO����7���`�?��ȮT�X,��U޵�8��w�������� ����)xg�Pk'���;�`޸.40[}�����vwS��
��R:`����$G�!m\���|��-�~�e���<�DA k�p�ۛ��B Y~B�-u������Ĉ�mB}as�Viy'��-�:"���ٶ��`������e�5G^�19[��|U�X	��ZM����k�/<x���OC�`���.�C���ɠ]u��Y���ڄ�$,ic�Ls�Ɓ�T�:�'��c�u4���Pb/��d��?f�|�����򞀱��[�\m5����^�̕�*Cz��C<�#ÿ	<�`��z���;(���4� �<��3zG��Ɨ� 7�|i	5� @7n&pA0b���6r�J�S�~9]�sԯ�Nt$���J!�r=M��}��?�*o���.O�=q���x�jV=`{�xR,��'Z���	���n+�,����'��f�w��e�-:-r'�Wr��t��+��٥�pS�#�\�@���0����H�;�����VU�	��*v�I�I���4$�����P�^�:{~��Q�'�{�0
��1Ey��Qʈ:#����3��n�{��J>_�rh�nU��?�D��G��pV��r��ОR�(v�J�=��E)0�`�GiJl_�D�`%���cp��+R��b��5�j>�ߨ�l
��*!���(r�o��r��҃�x$�_����p����Ab��1
�
�)���ad�Ea��%-���S��(���$�O�9%���@�"��G8ki_�����wn����@�ݘ�ícM���9s�NG���Ec�.��.(k��%Lz��sp��qX�A	��.��a{՛D*�����cB���7���F�;,1��e�4��g���Q:"Wd�@�89��R	�O���R
����J�>~�.�����?kd,k�0E�!{4�-0l��8��[>_6�e�m��q������y��n�y0��Vgy��ӣ#@��`4Do��D�e���1�Bg�nit�p�INS����3��6�$�j.�Kq��⸖�Y(�G�K/���aT��K
3�5-5��3�jZQ���y�]Ein�_� ?2r���D�h�����m�����/87Y��"f���g��{@r�ƐT��KΒ�.���ξ�����M�őB�es2�~��0�*����d;��y/��e	öUt�>������1h�G�-��h_6�b��Q��k�a���!qȇ#\�=�N�O�r� �WWa�6���[��5"�����'��wfA�M�W�ڙ�f�S~�tN�r���ٜ�S'u.m���qӊ���(�P�O�ke>w@��,�?!�!�p~�ҙn�R�%*�%,GK���2��S��\��u9�#¢m�|�R?�IF�R"pB�FO,NT��E"���r6�xr��<FO&Rm��9��@H~����y珬g��|l|��ً;Tu����La�5��)���S?�����P���5z$��Q0>�����Rg�%�o���8��o��=B|�=�� �(��w��8c������e<���t�,��m�A=��@#�6��&x 'J�9����-�*h76��HQ�\��(mh�	�*r71EV�n��ֶ=wwe�4.*�şV��[2j��r� v+d��yY�`���6�Zv�s�6t�א�K��Nڽ��R{�\;�_�*�ѕ}T��n�T4�k�Lc�x�rQo�9+�2c�V��״�]�_�5x�{�f(v���lum��A�gE�5�vS*V�(�<&��_0��QJ��S�~A ��ye� �Ǒ�.ː^�ǩ��ˏw�{�詸i*2�m�����G�X���9�#���O�eH��gs
����}���_A/M�1'�l�	� a������O����(K� ��b��Gxl��Z���h4ԓAyf����^��P4��b�>	A#_c`Z6�:��-j���Xo����ݪ������Ԧ��������a��B��{?[ퟏ������Q_Z�4d������h�b�|�o��w"'՞������/�� (0 ��rr��f�.��ˆ�;�����"|��{zð��}��1��a�TU�J�͎(p�o�["Y@�f���)/�cY��.������P�V�!O��UD��u��$��1�%}d��C]��	���@"M;�ިU��'S=ʖ�t�_9+�5#*����3Xx�2H��){����K����*�g?y�Q��y�����r��h��+��B���|~�.�@㨐��ٳa��0*��!ܺd($�2����n�v�}<�.��B�7�/z��l����t<� �+_��Y�IZMB�	��xt{P�T���֒�HB�f0<���'�q��+�-��po�C�E8a�k�^L5��"9���,!��8����(&�9"t��Z�\KT��:
�O���Dz�Bi(��4�/��X���Wm�<�'y��V�2����	��%eX�����F��:�c|".�5�6�(�0t��B}�jff@ʲ���ɹ�Ű�u��^p�������zs�E�=�?��:	�R�@�zL�8�5I��hdA��v%^��A`���B��!'�NA�^��������枅�y��H�-�6�c"�t:S5� <����6�2��䭪v{R�������Ms��	�S�"˙�O��R�7�T7�{�_w��y�2KNȢ}�ᓇ�CȐ��칵b����>���x;诪�?��e��C'݄�(Qr��Ɓ{ '$o�~�tN�P��Ѐ����D7"���,�Cz����ߍSQ�-��+�d���µǼm�Yډ�y1�%^����4�MZ����f���5��Y$�:?�zHi��ww(��%͚<�s����h����７�A�)�-HY�t�傘��+f$*��u�f���='r�,<Y-��"�AC�&��-���|�7���-�R�}�0��m����|�cO?�!�]b��f�7|��m�~�9A���P��(Q3�3�s�C��W����c���$Ik,�IĘG6S���$3�^��`�!v���V�<c{��U��(y�=��[��Z4@�L ߐ����yP\p9���U��*⨢��&���)��
q�l]G��`ne����D��	�aT�M�vǥ�y�Y�N���K�zC� �q ��u��P則U�k�#�}������o�u�����l�)<�H�d2?��+�	��5�Ɣj��
�O�􏄾��1���#?���-�<�/���1n�!�w���� 7�Ċa��fG��[��6��1�� Ɨ�W}�e�AOB���P�jG����/���_r�J��'8��x��|y���P���>um�h� D���Rj�*P��?�
���X��@���n��D��m�Z{-j��~)�'T��ru{�R����U�S��v6�-�f�Kk�k��!�Mvo�&�,Eߑ�"N ��N�6��f1mT%�� 0�ϯ�:?E�r{yEw6�@օ���v�M2�2>���<�07���8K�ח��{$���L��H�ز�^HU$���7�%�嗀ϰ�t�z+����H$��r'2L��pP�ny�S~�ǃ"��Q�9��&��\ �⒥����E��fDrWW0��f��|�F ��C�ݺ9�����͆H^"�[n��M�K;� �l"�[��\0�c�3�\�2*1:���{��!:���d ��Rm�څ�E��I�%#���h`�J��Q�����l���P)@��Z�°_��IS��R�o��?�i8���l.2T��U(3�Y�̟���"��{}��L�R�����\j��~b>
�rb���$ռG$��y�q6�O1nԝ�\��!n�.���ŀڟ4^��H��	"��&S�*�
6xF=��3
��2n>i���%� �1�!���|K�
3�rQ#�d��3h2(�����&p�d+���hJK�w�������t��HG̹p@,͙����I�+m��ՃOյ�w��6�Zy�J�Z����#���oj��a%]Adp�E��2Ѡ���Ւ�[ӑ����R0N&_��v]1����+$�^��_;�r���Pi����L��f).:���^���^�Z����#~��g�(���h�s(�;��̤�IyZ��
�O��Wȧ�A�B����,=�S��)��ڛ�Ԏ�yV]���$0�lj�7�<#\"i��~�7����6!�_G,���G��f�k�2K����-�b�~����ʃ����u.�7��(Y$�(�_Z����:��p��8&��}!>hUIΡ���J����p�		=�q�]����{&��q��,�H���V�K�����!�\ɽ�#v��zʠ�!��3S�m��ѣ
����O��aNY�w�	����Ыل�<L4R�L�m���&d���j�A�γ�c�U'��^��M;� ����R\��3԰��Sd�o���e �_5~����zj{���Y���ܸŭ8����r��n蔹;y���[�)XG��V�7��bzRk����K���7��-"���|�s5���<D��_#�%��"ݽM���7�Nr~���1r����|�$��L'�u�~v`����vj̺��YmR���~�+��:�4N��Y����)��L�����w�`;��@�ܲ7U$E�a���G6��3�4�9z�ZYK��v�� ]4���}ږHbU���: �'=�Jn��P8���i.�s���k�pw]��t�!G���*`��ɲ� ��������fK��s�Ւ��]�J�aymX�^_�I @r d�b��q0�����$���o�~��B�b_Jm*6�őԐ1�M�y�E�6UW�ڧ��p� 5�{��Y��5��Pr�-æ�W�yL�zrP��>����S-l7ۆ���.k��E�h+���2�|��毞}���׭�h���8�Րf��6C]bm[��3?�`E�{d%!�6��"�H^����\{��l�����T��?��tR��_,�����Z��1� �"�WC~�H�Y/˿�X
0�(�L|*S1A-�]�ߤ}�tt�&���{�)5M��\Z��v�h�A����g�n��^�em	5ix�m�b����c�wU�h�%�!?�<i||I���-��Z�FAϳ�y�5Dj�Cc��txn������M��k��K�[yw2ѐ&]=�z~H���"���ޜC�$s�D�ē����C�Mj���Ơ�'����f(��:/Q@��DS'.��@�C�G"��W���(L,m��9&LT%v���IpYۿ�&�S+����'�y�2��Uo�*�Q�eT��%'.734|����&: �y[��}!4�����X�ҵ�x�#G��u����۴*ӳ����%���*YN���BӮ�7ɊN����E��p2��+�/L�g�&o�!nK:Ԟ�Np18���K�'kI�8��{W�� �PP0����e�&}A�"9g�W�Z9[��Ѳհ��~vo�2�%��9�э��ay?��o�a�{�)GԈ��J��R�1��8Ή34�6 ��]��<�n\���A�y�UgQ�;9
�����&�[�S4\�R��D�ٽC�-GY������b��Np��0V�;q��6+ϪC��uT�J�H[w@�v��n���Q���T�T�'��k�M20405!o(���Sev�;6�cǊk���x�|�A������<'�>�שu��D�t�d���~n����\�����'�a�����'�ˡ�X4Y��\�����������w�nmP���ћ�3.§)�L��|C��܉�A��.7U��l�{o*��	��B�I�_�,E5�R4��΢���b��,�%D\,��}aҪ�j{% ���S9���EP��������`�&/���W}��Fżv/a�i�k�_S_2�.�����Po�\��S���*�g�C�\m�w�rK�}]ħ��ɛ�h}�R�I��������K�3X#̣��r�����ܓ]��;n�7��9H�p���q�?�Vuۜ��uF~��'�29ݎ���S��$�+���c-���vId�ڵ�O�@b�V�u`����bڎw}A��Q��LƎj[��:L~��Kn�.��;��$��=�/A�^̸�X_�H۵���d��\�.�Q̐RY���p�c�3���,�uPQޡ��~e��:�}�jy0p���Gtţ��&+ȓ?c�G�l�+B��:Ɏ��%�&�	�����]����~�/+�Z:E�^N7�U~|��s�yI{���\30��}�uɻ1@|��0��Ю�w����e/�#~=}��������-���p�it���w�������]���"�C�P��H^ ��:_m�\�9)܂I�/z�D?*�)�$:��0T�õ�C4��;O,`���:|�!���uH5����Q�0@����F������.�%�T�(��')�}	��}���~B�!�] ���ET��[gV7,8��;�H���h���|��1�����#�MZ���78Y�q&x�ib1Ͳ_}>�8�A�H�/�)�T�1q`ewo�n����b!��Xت{��RG��_v�/��Xʲ?(�貢k�I�	;D�a�#�i�)����C1��S��%:��֔�9�����k���0{ݫ����'^��GLXL��P���s?}9f(����[{*[�Q���Kzr�����x6�C�����3n�K�T�C��P��1\F`������$�Q{nŷE���� ��μ
��Gju�tК����<Mȑ%�P�yP��#�M0~�b=�����׭��׸2Kb�5��Q���B��yA.���Eď�r�f��
��M��ަi�q)=i�*�݀��*,��u";��2t'�a$�j�P��k,�^�a�aB*��Q�h$p�P��ᓶ�����T�p����m����L�M��ѷ�[`���-�E�����QXļ�X������V��!r��ٽ+o���l\�Z�����v���7"T��-�F�#�w������x�6Q���
1�&�{�뺥"�%lD�����G
���͂O�����{��X��B�E!�l�\�0	I��ElWz�=f�]�4�S$�s�?ԕ��?i(F����؇�����쒏�M�Ư�����;�5b<�~%�,5���S��PCF(=R���Y�N�tsǡ4��q۠V/��r�ٚEE*�W'�b�x�Zc�\�L���j�a�E�EЄ�k�k��ܳoH�@��gNP��&AQW$�����Z"�YFX���B���n��\U�^٦����½vL����n��&�$�ϻ�6J�3v�������Zw��_�`�j�;c�a����#�Q����������TE�	�ir
w����JZWg׻_Ʒo���5���L�~�u؆NZC� �D/J%ګ��� �dه8u�Z1�Hz���4�m�o-�1�B�@��}u�����N(z�Z��ù(�҈��#Vo��%"r8<S���Z�`d�S��)HI$y�M'��+\�[��yT�?�0W��>��A�8C�������p�W�W�N�|��:x6,0"j0���.�KIx��!�<5�ͱMӕ7���g�l?��Zfe3�j�6)O�k��&�� ��5����`���Β'A-�g澒�^e�SGGX�����W4",��(�����c1�s�=p��(�VQt�(NL�{�$�$�zW���./r%ٰ��	�#p��s�m��Z%�~�i�}��9�%��bj����ߢ�c�+V���_'��7�N�d�秪�nmz���ٽ&:��`�m�W��Y;բ� a���!�M~F	ƢZ��|2�.-�C]ؚ
���ŋEj��2)�Ck��@#�W	�V9��&����^�%P��LM�)0�|1��AP����>N�2d�ٶ��'}����v�*��BARO��aZ�f;�r���"G���=B�P�*���$p
)!�9�����
�Č��|Hö���Mj�l�� ��$>�ʽ^�ޞ�����{��E�2�J�w�DB���7&�>�j�X�R�؂��20:�ylѴ"�!��{CT:E�c6�/N^m6Mq�����xƭ@����
�|7ĳWG~	A=M�j���a��������T�)7��'��7���	>x����M�nL:��/��+�'�>%G6����9H�؃���3�Q/��ie�D����3ɢk�ߋ^�I�ǩ���P*�M/���i�g	O�q_·͊�o��)�����j�Z|H�~�tĭ{��W�"���"prOc�~�b/W��'_��{��Z��w�!��$�G�O9�a����Aÿ���s�^мNy����u�hM�|ee�WH�Br�|iҺ`��@�eӹ�0�ak-xL+�"J���И*(��R�pL� )H�r.jlf�_�OY� @�y�t�I3f�豅z������0=�y$��ToE��N�t���d����
���N-��h��J�9�Y����;��#U,�����������%f�⃤�c��%@��;��bd0���O�k�C)ސ.�	��g��oޒ}e�n��]�d.N���H.�󲆓�u��fk}H>�,�a�x����*;HU�<���+Ð#쿫X�;����?��ćLh��ŉηH��#e	r���x�o��[{3�#P*�o�'�,���r�2<2q���xc� =~���O��;O�͚� �����ɎV�;l=-g���5��2�����yЄ�8��g�Ee���=kc�Y�>{��O��:�	4\\���&��
�J�X�J"?�H���n:��4���""�$iW���FU�g�e��x
e���79�a�)�)GY�Е��9�f�����~��]���jcH>*����C��%��.�����"Z�m�O��O�5f YJb����gc>̨}�D�[��ۗ̏+Q��E�\P���oq�. �R�mr)�
��n"��pL4����CF��� 4l���X%�� K���+YVD��6D[43'ASpy����6gQݾ�c�˪�.��W�Hae� #��\�:=�8(��(5h#��s�$=X} O�?�2u���38�Ϲg����@�<Ŀ��i�� wTk@[�����B9\\��+[���e�Z�rxS�T�!�h6��֯�/'��	鋷n�j�\.�)�&Q���,���xU-(�ڧ- bD�cy&ٝ�GDEEt�� �Duԇ?�~kW�kB������� -�(z��� 6z��q6�I^��
�DU�3E�����1��#<ej���XD��ė��q|?������q!�C�)�vT1�a�g~Y=��TA�Y�PP�dAs3��5=0�F!x���[ɀapͣ�t$�5`
as7	���6�]�y��?�'+V���ߘ"$�c�]/6:7zJh%�Z�m��l���,{�j�Z�es�s�k<�y�n�fz��x���]�,^[��u�
��}�C��#�8���k���R�c`��N�Hmm�02jU���w�ֱ�jX}�%Q'rJ������� ��֛���s� ���a�� F1�E�J��d�AX���g*�/��)~E��Jձm]��ai�U�|{q���h��E1�~'�_�W������4�G!(���Zܒ�l-����H0�(�҈o��(�P
j����蒒5�EQ�-�hz_�_�����n(�d[�[RS�e|�$u�w�U	�8ы�Wk�?��NbQ��`��F����nCtF"�	'hA���l���W�F�3� �����2w��^��LL���b�s¤���8��
�w�� ��vz�Q�n��G_�]3�G�@�v���)��pm�C�.���$�}zMA��d�ZH�FR|�h6�X(����`��U���0-���|*02�l�b�mΐ�X�����-����gC�7�����O������1��	T(�<\06����2��ϗ�L��\a�M�X"#@�ۗd���]���L^��H�2Y\U�8S1�'xq`	���BwL�tbh�ra�%�4Ė���j\*�ʋ��xX���)}��~����W����Ynd�E�U?�kZ�m7����(�Ȝ����;���I���L�E$���ײ_֜�U���).,�7��cAf���CX]��>N�x�V�r{U��W����:��4�3}n`A�:�#y�h D?f�ǒFY !a�p��+��i �幠��f�۱��o�l���ٹ�)M�2�^	���sM�(��j�<Myi�2�,#/-�q$ƹ���� .�ö��B6go�B�������f�V(e��ř�H��6�bC7��2e�ǏTT�qp׼g�HtL V�Ҫ<e�a���4��IYL.G����Y:�Z�F5������W<� E$�Z�v_6����& ��=��?MfI���R	����1Rl��k*<;��������9��P��6̕.�LT}8���^p'���@��-�Z[�6�՞��A/��6K�55N#5  ����Må��F͐I#�&�V�R�m�]��@�"��t�?���L��E�#�pe�������}��7�W,����+�ETh*.+G��%"?{�<y�$��^���ڑ�N���F����;x���)���~���*�F��SBX7꜈-_��V[�Wq�4{n���6�6U{�P
�o�͊˄�&unM���R�9ѥ]�t���kS�vMZX��L-�<ӹtK �nĂf�<����eW	����u�Q&W�W����w'3��*=ZK��]	�7V��g�/���L�LcnH��1iv�f�{����ٯN��d��LR@�vim
�������V R�ٚ� ]?,�`�ZѮ��H�n�\p�,p&�f��P�(76m_�|�LRy�>w�Ī���]?ן[�f*�� �W@ᑳ�M1��*��҆���C��/�hg0!�jT��b8G�b�%	}�e������ZFh%�l�~�~�������s�΅ ��[7��m;�`ܙ2n��H�O	f�����σ�Ǒ"�%c�-	r���%Wz�RNq~�C 8n2��[���|Z�xk��6}�M:h`��\���#�2�8�B&�12�ψ��}A~�L�e��k��k���y��p���y�����!5��g[`v]A���ٕOQZ���|`G���7�餝���g�;�޷��`/�Yǝ<s�����˨��s.Ȝ�>�\,�iE���ؼ�o�An�|`����L��!� *�fXB���6@������Z��]��D������1T/�Y ȗ2�spg�M���kw$M�{�`�Dݼm��P��H�1.�Bӄ1����������;�}����l�h� [G�&�2o�B:�����W@j`�w��~�Z����B�]f" V݈d &���e��W��ƛ�lc,�?��X^�+�JZ �cg"�?q����#Ǹ�6�||�|U%�W�Qev��t�ػ7�� ����,�S����&�!�I�E? n=�m�^�P��[ ������)�a8K&٨��g~�A��
rX)��^���m�ӗ	�§m��Rw~�k����L��D������C�@��bo�	I>����h#B��#P=ib7�}�x�R��5,>X4t]t�jQ��5Gl��� d���]q���b���AسyۗW�h
��k��q�X��[��|���4�<*	���D���.�n�)+z jb�
r��v�D��
�QY���e��d��s'�G��;X!2q.��K���r <��,��Ӑ��@��&�`CE���|*:aLoOTvu���P��.3H�/?.D^��9����W�`�
��2h�"�9U���h;��m���9�':Ð�m�k�#zd�u���ܐGS}���C|L/��'�8�'�?�x2�$c��0{y��K����P���>b��7K#ʽ��J��8�#;���v����YԔ >�iS ���k�'�z#�p��D���gώr��%a�O{�X���I�a���K��߽��I��Y�c�V�U3�u���)�_/^�J���M��i�/ۣJ�2��k�R�}N��'��ƶw[2�҆�J�R�-Ve�.��-B�+�#��J�hP"E ��Mz5�IW�W1MlE}3�V���I(�R���?��Y]@�P�5�A�Fz��>�i�+�MXӻ�r����.f�<�pFP+!D~��u��WJh��0(@#��-HV�VҎQ��۹,���Q�=��ٛ�6駍��b��"j��j:��U��#x��wk{��W¸�G��}B����Q��r��\ϔ�ʇ�:N@�[=�O$5ҽ���y�I�:[��kK���C
qM�<�'���X+0i���#bHf��̽����c!|�ㆀos���^5�]�0&N�I�|M�Z���ͥ��Ű����W�\|��Ap��3B:�xN	A����?Z��b�*n�5g��u׼� ;�m#&������t"��!��z����絏S�4v������d��LF�Jd��}]^(X@�Y���U�Ɗ_�L��,X��籾+���rV���&㉫�ȧ�;</�p��%���.`<��e���+�F�Ͷ"?����
�%�B�k�;à%ᗭJt�%m �;�R[6��`-��p?������	�,.��"���"{�?e:��
������R��V�X�~�K��Gp_������n�!-�dD.�:r�i\2�)����
��;�
٪��� ���Ҧ�������3��Mv9q�D#[��I''�'�J�O�"G�5p�eL��%������qO��kH
�X��V6��xo:���%�=ok=��C�/C\!�xV�w��NF �MrmB��|6��yA��	���j��9*�8�d{P��D�F�"W�VJ��q&�j�kz�ٔ�r��v����K�(E�i�@֘�o���Q���e*�[���(djE��:HsWk`��=4Pj�UR���[߷z^и^��ݏ�C��e���7�9�7zP���Pm ������C<�{�0npș�e��of�KHJ4ќ�C�jL-����hm% B/a�ϧ���VL�k���Lxt�q���|ձ������F`|;Dw���;��l���f�ȑ@e:���Rc�P�lG�?챦��(��_�ˈg�g�1�i#�_�+��6y�/�p@���/Éa��ypi��w��|{���C�*���t[�;��wN�V8P��hMh�B���P��0�e
u9����6/�}�#���C�6A�g|@�Yu;S���J.��{�׹�� �G���� �F����\a��V�Idu��G�v��3&X���.��+O�����*�N@�uv������Z�Sq�����O�{�cnZ�&��l�d�D^~��G՘��v#@`ĊISK�`�2��[�I��� �rny7�!@������W �Ly�/C4������|
���q�c��n� }�I�nQ8�E�k�>/>�����z��6KX���˝���x]�x�w����AM��i�_���*ˑ䆒�F�����d�:�|�d��4�������KI��y�<�*�ܩ�r��@#��)kZ���j��aJ[Z�9}4��A7��ul_Vd��T�~0��/#3�ݧ-فz��Vl� ���2�R�9�aP/����,�RbM&e�^lĦ=�r�H���Kr0�@oC�^O���ͽCO�׌�C�ɩ<N��F���`*D�����x�*���[����S����u?0��U������H��^]^<�4!�&�O x/�>�@<ΐʧ��n�?��4���𾪰����Bl.�[h�y���?��&eчX2YY�H�L߷�H�j���"D�l���z�w���r^r�̹�Fã7�)������1�ot���'<r
��<^Ҟ��.�[�T �n�
�K�V����]^/,�¹F��|�y���>������ү�X%#�b4����?����0�GUc��;��'G���Xj7s��><��|��:�:.-U!�&`�M�F}�ݥB�~��t��t>�!0)�w���*��!=�E=cQb�uhL`%ữT?�Ts�]�*$n����ڇB�D��.�����������e���S�C�n�6j�UJ��Q�!i�5�Y�yW��} �vB�mK��f��D�W�,�6 ��� s��������y�Z%��U�Ө$�$d�$�2�Y�%����,[��j�r<M%�qsJ�=K��xˏ>�����+��A����H"j#�8[����+�
!�nx�T��@AĄ㌠IRA[��{"���"�	�!^;�d^-|K�ݔV����^�B�p@YE3@�Guӗw������>ڟ�ih�"k6��hӣ�S���#�e���Q$���Q�tp2�lR�/DR
�"'_���K���ٍ�^����5�@�V~�*=��y(�ݫ�^y�� $�y��N����;>^�f�鰃��KLl08@"���[�n�K�����3*���w�~�qe��<���b���A����x�u�۵�ؚ�J]��s�0����2yE��������z���]�8���$ҭ-O����
@,�0��V��|�U`�Gp��厷��tf�C��P����-"r�
<+��(�-�¸���q�Bӆ�/Z^�	�:�:<
������/�Rݘ��ގϳ�8x���7_�?Ź�\0�UgJg`Y��Jt��Q�+2{��Hm�O�[&��}�d�%���25K��yN����He�?m�%_�e!����d:k�^	�d���$�ʱ�����AO�q��:,��5�[�w���`��_�ں������2;��]��<�j�J�=��n���|@��a�(=	��gS��f|���q�V��`n<+Ʌ�CA�D:��#!%�V�{��	�ixÿ-iv�Kj�첹t��[x~ż�s�=��R��E�`���'�N2$_���]z���/	A�5r㍭g�����*E��F�#�}:̸�|����>��r�44!c��]�(X�筿xl|I���Ba���L�l�`�;��z�+�ٷ@u� r~9\.S�g�:����=�%ti���_��y\�3I��*�JH;�b^Q��2��\c:q*��7 �5�Q8�R#O͖ü��VPB�BpO���\.�nk8�j*X�H	_��]�� 	�6*a]�Y��#*�+�NH43�/�����n��i�\���0�v����ښ�2�,P6I	_�o&�wk�y���'&n�j�<"�To;����S��[
�Y	?4��"� p�4L �ԌYg/'��C�6�`t�"[.���O��y�0���/���W�>����T�g'��b���"�9�$�Ԭi$��%Ηȡ��yӐ.��cXW�\EK�:�c�$�'P�w�8w�n*h�-���Y�)�g1{u��%�s���,C-1����ةo$���
�"a�]m��b�̮��z� Y( �͓��K-�r?X�6��L6�7oA�Ա�N���D�\��R'�jص*� ��YՔ +����
�e-����)�]6�l4��W����I��'�,ĥ�Jv�t)��.�i�gU��M��
����i&��r0��Z^��6���yv۱F�/'5e��`��(��Y�'�ʬ;�����Gt����P+gU��4��2���>`�H�Su�˄%D93�D��f�|���6$P��;��hI�rK�S���{Q&�h���kN�lچQ+��Wn8��`މ�`5�k��61�d}�"t:����׊���9��l_��h�Y��<�␫��9��9+�E��g#���/�k~4����5#.q[�[�-��^g6�϶i���X.�>�/�t�\J]��x�6IAW+���I��IW1��kV�w�=�n���z����'��HG� ��䦚Ǻ�Lr���"#�`��5�֣`�ѥ<e�^;�gI���&�Qqp�U��5S�Z��:v�3� �z�5��sE� �ڥ��<�UT�dzF��;#Qj�G�i�rU����F���1�l,��M�I�"z��b���|)}]�{��U����SAj�1���}#`��8��1¥���1�j��q�Y�{6���N-%�f�#a������w�u#��b�Q�(p������l�o��7����P���&�[}��cJ�.�a���<����JWЅ]��ryyr4Z
��?�(� :��rR���8���Wi��.���n��H7�*���Эi�ɂ��}�=�0�Y�U�3gD�8쫵�G�md�a�I"<���0�^�c5�_�*L!��+}��N���\�APjZ��j�o<�"��r}g;�7(ma��)R+�i��U������|���72f!'u,��@�ٚ�a�O:Լ�t���>�~5"��F�"X��&�{�q���}�д+]�tB����w�j�ii�-��gy��ԟ�3���V[Q���-�B�z{tq"c��r�̀X�/���A���K��)a3L�l����3��-��E�K;�{=��.�ا7CЎ����
q�k�aa�/�W�jO4J�-�)J�����-Dq�#E��HR�֓�q%��{Lr���ֱ[��~H�E�O�$zȳ>��p!G�yr��·�V0�Me�d4B�Y4:���UtqN̈[���:���4,��A�~|@�*4��(�Xg=��x���O4��W���	q8@��D���N�.���|�yq���<�q��[�o�&�J�b��MR�`z5��%�߂(m����hg�}���Q�k&o��m�t��p>M�o���Җ�#�;oإ�=�
H1�Z6��N��E�"~�1��~Us���;�dq� �3�;zD��JG�@H4���Aӂ��0傰�nf`_A��d��[TkvO0�Z����^�jo�5\��l��4���CX�`۫Z���S<�g���9	�ޑ���
ED��:D�(;W�nݦ:���12�f��N3��p�(�	�v��)�#!��.��4-V���k~/�	ye�t<T!��̧���\|�W�Ly{�GĘuv��z$'D��WAmpd�<Jc	�8�|5��+��0�Kȸ����Ǥ�J�:��I�ś�&%ʐ
N@��ޘ�n����WUY�Ω�]��d��I��di�}�J$��C�D�Bh��\^ ��U�����V���h���F�* �6�&�DL΁��S�7��@�5���A�����*��8 �Rv�oő>�y��C��w�b���f�{K
i��9�1m�3F�c.�lPn�����QN9й@�O{.�����B��M�`�����&)ɍ�'㺧$Ǭ����A�J��(/��IL�l���7�:���Z����3��רN���j�#��fw$f���8$F�ݎ�bG��$#��'�1���ڏM�슺	�O�k�>Y�1}�@Op�ހ5�����1�d���l�&
}�.r�.}#����
�*?Ϯ�S���iK �ͼo��.�{BQ��K=�v�%��h�ҫ伐�� �jF�4(x	�D�����v�D�m��#l6��fc�9<s_[��J��<��2�
�W^ʖv�o�m��=�JR�>?L�͋7�{��v�!6��ȱ�ە Dx�1r (߉�I*��Tϭb�f�J?��fA��*D�?����W����`U'�t[4�u�bAأ;�Z���5��*K�`[yMU�S�t��rj� ^sB��B�����?��L� ������L��G��L��:��MW�� E�T�M�`rks�6���no
׎�㷽�*�Cn
����"5���x1Jw�@;�e��ڙ�ŭ��fᥡtՆG��5Ip��Ki��
�X�]bf���>��&U�ݕj���F/)�h������ܳ϶���Æ�QV�P&���4����������Szi�Q
c���9>]x���䝇�����Պ�U]7?��S�Z!�IUjAj�F＿�vīuP�ëNu��!y�A;Û���!�`4XH��3�P��S���n��,�'�V=�l'�/+�ĺ�zf���KP+��\�9�3ȧTvA����"������4���*ڸ���S��EE�����(�<�^Ns}�L^�!���y�͍{.6�h�%�2�)�N|4���̺����϶U�O�y�8�%Q��BY/L��'�$֘�C��c���C%�� z�Ϩ��:�J�.,[��}�yשUL��X�b�26���*���i�z7˫v��l��CX߂�Ʌl��[�U-�[�aNd*+S4��z0?o�w�1�3}�䅲0�o�)�5��J�}��Xk =��Z�B�*E`�V��C�W�e��#�J�������C>Z��2I24�������=`��[.|�n$X�����v�-�����=�1K��Et��6:Qßo�M-ygϰȧn�	��M�`(3��s�J_�� �O]���q�n�+R.\��� �*�H^m�̓O^��S�a�9Lu�-�W�+�GAoiQ%xJ��oL&�;-�?����\$�&:U��kYr?���h)�3/�Lv�`>ge��uP�;���c��������E�^To��ӏ��}�$7*%�y�|?�n	�q#�����>Q7�31~���0����,����'�����W�
���ً�\·8�b�ʗ���V�A����2rEP��p���!�=ՐS� ��>L���w%��ث	;���Ȍ���ι��`�2�������F�)R�j'�8�D@~e�Ԛ��jY���c�Y����Jd`�x)~v%Ő�@�c�?�S��R,K*mk
��R �0G�E���n�#A�&U��sji�0м�S��uȽ܉z��I���>	���v%�m2y{�s��P6^�k��n�>^uG�_2۰o�"��0����w����n���� �G�=��7���旅g8Rv�ȱ+��
|��?=e#7|�F0�����ت8㈄� ,=5L�b$}�}K$lp�e�H�ۘ�={
��&�گc�qO����1t�<�[1��T:#�5A�� d$�]$��~0 ��� @h,�f����^� 	ӱ î$z�Aa�9�ǈ��A�3��L?b`9=&����{����;�g��K<�2֒�վ/lu`ծ>Fy^E�[a[ǯV�v��B�һLRtX�1�
�u�G\�m��b�63R�|�-�_��O�$a������k�hn��_���%�?��$5�b���8>���%����7�S�5����g��`8�+l0B6Қ\�U�^���_��ݑF�>Le?������?ժ�l����<,���S���V&}���祴��=B������ �S�� �Q�a�5�G�9eN����Z�j���(�D��]'V�<�}0unB��Q�=Wt�k���9#0�8|��4RL����e���j T�V�G�yu#���e